magic
tech sky130A
timestamp 1702613480
<< nwell >>
rect -70 190 1070 330
<< nmos >>
rect -120 0 -105 100
rect 25 0 40 100
rect 65 0 80 100
rect 130 0 145 100
rect 195 0 210 100
rect 340 0 355 100
rect 405 0 420 100
rect 470 0 485 100
rect 510 0 525 100
rect 575 0 590 100
rect 790 0 805 100
rect 855 0 870 100
rect 920 0 935 100
rect 960 0 975 100
rect 1105 0 1120 100
<< pmos >>
rect 0 210 15 310
rect 65 210 80 310
rect 130 210 145 310
rect 195 210 210 310
rect 340 210 355 310
rect 405 210 420 310
rect 470 210 485 310
rect 510 210 525 310
rect 575 210 590 310
rect 790 210 805 310
rect 855 210 870 310
rect 920 210 935 310
rect 985 210 1000 310
<< ndiff >>
rect -170 85 -120 100
rect -170 15 -155 85
rect -135 15 -120 85
rect -170 0 -120 15
rect -105 85 -55 100
rect -105 15 -90 85
rect -70 15 -55 85
rect -105 0 -55 15
rect -25 85 25 100
rect -25 15 -10 85
rect 10 15 25 85
rect -25 0 25 15
rect 40 0 65 100
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
rect 145 0 195 100
rect 210 85 260 100
rect 210 15 225 85
rect 245 15 260 85
rect 210 0 260 15
rect 290 85 340 100
rect 290 15 305 85
rect 325 15 340 85
rect 290 0 340 15
rect 355 0 405 100
rect 420 85 470 100
rect 420 15 435 85
rect 455 15 470 85
rect 420 0 470 15
rect 485 0 510 100
rect 525 85 575 100
rect 525 15 540 85
rect 560 15 575 85
rect 525 0 575 15
rect 590 85 640 100
rect 590 15 605 85
rect 625 15 640 85
rect 590 0 640 15
rect 740 85 790 100
rect 740 15 755 85
rect 775 15 790 85
rect 740 0 790 15
rect 805 0 855 100
rect 870 85 920 100
rect 870 15 885 85
rect 905 15 920 85
rect 870 0 920 15
rect 935 0 960 100
rect 975 85 1025 100
rect 975 15 990 85
rect 1010 15 1025 85
rect 975 0 1025 15
rect 1055 85 1105 100
rect 1055 15 1070 85
rect 1090 15 1105 85
rect 1055 0 1105 15
rect 1120 85 1170 100
rect 1120 15 1135 85
rect 1155 15 1170 85
rect 1120 0 1170 15
<< pdiff >>
rect -50 295 0 310
rect -50 225 -35 295
rect -15 225 0 295
rect -50 210 0 225
rect 15 295 65 310
rect 15 225 30 295
rect 50 225 65 295
rect 15 210 65 225
rect 80 295 130 310
rect 80 225 95 295
rect 115 225 130 295
rect 80 210 130 225
rect 145 295 195 310
rect 145 225 160 295
rect 180 225 195 295
rect 145 210 195 225
rect 210 295 260 310
rect 210 225 225 295
rect 245 225 260 295
rect 210 210 260 225
rect 290 295 340 310
rect 290 225 305 295
rect 325 225 340 295
rect 290 210 340 225
rect 355 210 405 310
rect 420 295 470 310
rect 420 225 435 295
rect 455 225 470 295
rect 420 210 470 225
rect 485 210 510 310
rect 525 295 575 310
rect 525 225 540 295
rect 560 225 575 295
rect 525 210 575 225
rect 590 295 640 310
rect 590 225 605 295
rect 625 225 640 295
rect 590 210 640 225
rect 740 295 790 310
rect 740 225 755 295
rect 775 225 790 295
rect 740 210 790 225
rect 805 295 855 310
rect 805 225 820 295
rect 840 225 855 295
rect 805 210 855 225
rect 870 295 920 310
rect 870 225 885 295
rect 905 225 920 295
rect 870 210 920 225
rect 935 295 985 310
rect 935 225 950 295
rect 970 225 985 295
rect 935 210 985 225
rect 1000 295 1050 310
rect 1000 225 1015 295
rect 1035 225 1050 295
rect 1000 210 1050 225
<< ndiffc >>
rect -155 15 -135 85
rect -90 15 -70 85
rect -10 15 10 85
rect 95 15 115 85
rect 225 15 245 85
rect 305 15 325 85
rect 435 15 455 85
rect 540 15 560 85
rect 605 15 625 85
rect 755 15 775 85
rect 885 15 905 85
rect 990 15 1010 85
rect 1070 15 1090 85
rect 1135 15 1155 85
<< pdiffc >>
rect -35 225 -15 295
rect 30 225 50 295
rect 95 225 115 295
rect 160 225 180 295
rect 225 225 245 295
rect 305 225 325 295
rect 435 225 455 295
rect 540 225 560 295
rect 605 225 625 295
rect 755 225 775 295
rect 820 225 840 295
rect 885 225 905 295
rect 950 225 970 295
rect 1015 225 1035 295
<< psubdiff >>
rect 640 85 690 100
rect 640 15 655 85
rect 675 15 690 85
rect 640 0 690 15
<< nsubdiff >>
rect 640 295 690 310
rect 640 225 655 295
rect 675 225 690 295
rect 640 210 690 225
<< psubdiffcont >>
rect 655 15 675 85
<< nsubdiffcont >>
rect 655 225 675 295
<< poly >>
rect 300 430 565 445
rect 300 365 315 430
rect -120 350 315 365
rect 340 390 525 405
rect -120 100 -105 350
rect 0 310 15 325
rect 65 310 80 325
rect 130 310 145 325
rect 195 310 210 350
rect 340 310 355 390
rect 380 355 420 365
rect 380 335 390 355
rect 410 335 420 355
rect 380 325 420 335
rect 445 355 485 365
rect 445 335 455 355
rect 475 335 485 355
rect 445 325 485 335
rect 405 310 420 325
rect 470 310 485 325
rect 510 310 525 390
rect 550 365 565 430
rect 550 350 1120 365
rect 575 310 590 325
rect 790 310 805 350
rect 855 310 870 325
rect 920 310 935 325
rect 985 310 1000 325
rect 0 200 15 210
rect -15 185 15 200
rect -15 150 0 185
rect 65 165 80 210
rect -40 140 0 150
rect -40 120 -30 140
rect -10 120 0 140
rect -40 110 0 120
rect 25 150 80 165
rect 130 170 145 210
rect 195 195 210 210
rect 340 195 355 210
rect 275 170 315 180
rect 130 155 285 170
rect 25 100 40 150
rect 130 125 145 155
rect 275 150 285 155
rect 305 150 315 170
rect 275 140 315 150
rect 65 110 145 125
rect 65 100 80 110
rect 130 100 145 110
rect 195 100 210 115
rect 340 100 355 115
rect 405 100 420 210
rect 470 100 485 210
rect 510 195 525 210
rect 575 195 590 210
rect 790 195 805 210
rect 575 185 615 195
rect 575 165 585 185
rect 605 165 615 185
rect 575 155 615 165
rect 855 155 870 210
rect 510 100 525 115
rect 575 100 590 155
rect 685 145 870 155
rect 920 165 935 210
rect 985 200 1000 210
rect 985 185 1015 200
rect 920 150 975 165
rect 685 125 695 145
rect 715 140 870 145
rect 715 125 725 140
rect 685 115 725 125
rect 855 125 870 140
rect 790 100 805 115
rect 855 110 935 125
rect 855 100 870 110
rect 920 100 935 110
rect 960 100 975 150
rect 1000 150 1015 185
rect 1000 140 1040 150
rect 1000 120 1010 140
rect 1030 120 1040 140
rect 1000 110 1040 120
rect 1105 100 1120 350
rect -120 -15 -105 0
rect 25 -80 40 0
rect 65 -15 80 0
rect 130 -15 145 0
rect 65 -25 105 -15
rect 65 -45 75 -25
rect 95 -45 105 -25
rect 65 -55 105 -45
rect 195 -80 210 0
rect 340 -15 355 0
rect 405 -15 420 0
rect 470 -15 485 0
rect 315 -25 355 -15
rect 315 -45 325 -25
rect 345 -40 355 -25
rect 510 -40 525 0
rect 575 -15 590 0
rect 790 -40 805 0
rect 855 -15 870 0
rect 920 -15 935 0
rect 960 -40 975 0
rect 1105 -15 1120 0
rect 345 -45 525 -40
rect 315 -55 525 -45
rect 550 -55 975 -40
rect 550 -80 565 -55
rect 25 -95 565 -80
<< polycont >>
rect 390 335 410 355
rect 455 335 475 355
rect -30 120 -10 140
rect 285 150 305 170
rect 585 165 605 185
rect 695 125 715 145
rect 1010 120 1030 140
rect 75 -45 95 -25
rect 325 -45 345 -25
<< locali >>
rect 380 355 420 365
rect 380 335 390 355
rect 410 335 420 355
rect 380 325 420 335
rect 445 355 485 365
rect 445 335 455 355
rect 475 335 485 355
rect 445 325 485 335
rect 550 325 725 345
rect 550 305 570 325
rect -45 295 -5 305
rect -45 235 -35 295
rect -80 225 -35 235
rect -15 225 -5 295
rect -80 215 -5 225
rect 20 295 60 305
rect 20 225 30 295
rect 50 225 60 295
rect 20 215 60 225
rect 85 295 125 305
rect 85 225 95 295
rect 115 225 125 295
rect 85 215 125 225
rect 150 295 190 305
rect 150 225 160 295
rect 180 225 190 295
rect 150 215 190 225
rect 215 295 255 305
rect 215 225 225 295
rect 245 225 255 295
rect 215 215 255 225
rect 295 295 335 305
rect 295 225 305 295
rect 325 225 335 295
rect 295 215 335 225
rect 425 295 465 305
rect 425 225 435 295
rect 455 225 465 295
rect 425 215 465 225
rect 530 295 570 305
rect 530 225 540 295
rect 560 225 570 295
rect 530 215 570 225
rect 595 295 685 305
rect 595 225 605 295
rect 625 225 655 295
rect 675 225 685 295
rect 595 215 685 225
rect -80 95 -60 215
rect 85 150 105 215
rect -40 140 105 150
rect -40 120 -30 140
rect -10 130 105 140
rect -10 120 0 130
rect -40 110 0 120
rect -165 85 -125 95
rect -165 15 -155 85
rect -135 15 -125 85
rect -165 5 -125 15
rect -100 85 -60 95
rect -100 15 -90 85
rect -70 15 -60 85
rect -100 5 -60 15
rect -20 95 0 110
rect 215 95 235 215
rect 315 180 335 215
rect 275 175 335 180
rect 575 185 615 195
rect 575 175 585 185
rect 275 170 585 175
rect 275 150 285 170
rect 305 165 585 170
rect 605 165 615 185
rect 305 155 615 165
rect 705 155 725 325
rect 745 295 785 305
rect 745 225 755 295
rect 775 225 785 295
rect 745 215 785 225
rect 810 295 850 305
rect 810 225 820 295
rect 840 225 850 295
rect 810 215 850 225
rect 875 295 915 305
rect 875 225 885 295
rect 905 225 915 295
rect 875 215 915 225
rect 940 295 980 305
rect 940 225 950 295
rect 970 225 980 295
rect 940 215 980 225
rect 1005 295 1045 305
rect 1005 225 1015 295
rect 1035 235 1045 295
rect 1035 225 1080 235
rect 1005 215 1080 225
rect 305 150 335 155
rect 275 140 335 150
rect 315 95 335 140
rect 685 145 725 155
rect 685 135 695 145
rect 550 125 695 135
rect 715 125 725 145
rect 550 115 725 125
rect 550 95 570 115
rect 765 95 785 215
rect 895 150 915 215
rect 895 140 1040 150
rect 895 130 1010 140
rect 1000 120 1010 130
rect 1030 120 1040 140
rect 1000 110 1040 120
rect 1000 95 1020 110
rect -20 85 20 95
rect -20 15 -10 85
rect 10 15 20 85
rect -20 5 20 15
rect 85 85 125 95
rect 85 15 95 85
rect 115 15 125 85
rect 85 5 125 15
rect 215 85 255 95
rect 215 15 225 85
rect 245 15 255 85
rect 215 5 255 15
rect 295 85 335 95
rect 295 15 305 85
rect 325 15 335 85
rect 295 5 335 15
rect 425 85 465 95
rect 425 15 435 85
rect 455 15 465 85
rect 425 5 465 15
rect 530 85 570 95
rect 530 15 540 85
rect 560 15 570 85
rect 530 5 570 15
rect 595 85 685 95
rect 595 15 605 85
rect 625 15 655 85
rect 675 15 685 85
rect 595 5 685 15
rect 745 85 785 95
rect 745 15 755 85
rect 775 15 785 85
rect 745 5 785 15
rect 875 85 915 95
rect 875 15 885 85
rect 905 15 915 85
rect 875 5 915 15
rect 980 85 1020 95
rect 980 15 990 85
rect 1010 15 1020 85
rect 980 5 1020 15
rect 1060 95 1080 215
rect 1060 85 1100 95
rect 1060 15 1070 85
rect 1090 15 1100 85
rect 1060 5 1100 15
rect 1125 85 1165 95
rect 1125 15 1135 85
rect 1155 15 1165 85
rect 1125 5 1165 15
rect 65 -25 105 -15
rect 65 -45 75 -25
rect 95 -45 105 -25
rect 65 -55 105 -45
rect 315 -25 355 -15
rect 315 -45 325 -25
rect 345 -45 355 -25
rect 315 -55 355 -45
<< viali >>
rect 30 225 50 295
rect 160 225 180 295
rect 435 225 455 295
rect 605 225 625 295
rect 655 225 675 295
rect -155 15 -135 85
rect 820 225 840 295
rect 950 225 970 295
rect 95 15 115 85
rect 435 15 455 85
rect 605 15 625 85
rect 655 15 675 85
rect 885 15 905 85
rect 1135 15 1155 85
<< metal1 >>
rect 20 300 60 305
rect 20 220 25 300
rect 55 220 60 300
rect 20 215 60 220
rect 150 300 190 305
rect 150 220 155 300
rect 185 220 190 300
rect 150 215 190 220
rect 425 300 465 305
rect 425 220 430 300
rect 460 220 465 300
rect 425 215 465 220
rect 595 300 685 305
rect 595 220 600 300
rect 630 220 650 300
rect 680 220 685 300
rect 595 215 685 220
rect 810 300 850 305
rect 810 220 815 300
rect 845 220 850 300
rect 810 215 850 220
rect 940 300 980 305
rect 940 220 945 300
rect 975 220 980 300
rect 940 215 980 220
rect -165 90 -125 95
rect -165 10 -160 90
rect -130 10 -125 90
rect -165 5 -125 10
rect 85 90 125 95
rect 85 10 90 90
rect 120 10 125 90
rect 85 5 125 10
rect 425 90 465 95
rect 425 10 430 90
rect 460 10 465 90
rect 425 5 465 10
rect 595 90 685 95
rect 595 10 600 90
rect 630 10 650 90
rect 680 10 685 90
rect 595 5 685 10
rect 875 90 915 95
rect 875 10 880 90
rect 910 10 915 90
rect 875 5 915 10
rect 1125 90 1165 95
rect 1125 10 1130 90
rect 1160 10 1165 90
rect 1125 5 1165 10
<< via1 >>
rect 25 295 55 300
rect 25 225 30 295
rect 30 225 50 295
rect 50 225 55 295
rect 25 220 55 225
rect 155 295 185 300
rect 155 225 160 295
rect 160 225 180 295
rect 180 225 185 295
rect 155 220 185 225
rect 430 295 460 300
rect 430 225 435 295
rect 435 225 455 295
rect 455 225 460 295
rect 430 220 460 225
rect 600 295 630 300
rect 600 225 605 295
rect 605 225 625 295
rect 625 225 630 295
rect 600 220 630 225
rect 650 295 680 300
rect 650 225 655 295
rect 655 225 675 295
rect 675 225 680 295
rect 650 220 680 225
rect 815 295 845 300
rect 815 225 820 295
rect 820 225 840 295
rect 840 225 845 295
rect 815 220 845 225
rect 945 295 975 300
rect 945 225 950 295
rect 950 225 970 295
rect 970 225 975 295
rect 945 220 975 225
rect -160 85 -130 90
rect -160 15 -155 85
rect -155 15 -135 85
rect -135 15 -130 85
rect -160 10 -130 15
rect 90 85 120 90
rect 90 15 95 85
rect 95 15 115 85
rect 115 15 120 85
rect 90 10 120 15
rect 430 85 460 90
rect 430 15 435 85
rect 435 15 455 85
rect 455 15 460 85
rect 430 10 460 15
rect 600 85 630 90
rect 600 15 605 85
rect 605 15 625 85
rect 625 15 630 85
rect 600 10 630 15
rect 650 85 680 90
rect 650 15 655 85
rect 655 15 675 85
rect 675 15 680 85
rect 650 10 680 15
rect 880 85 910 90
rect 880 15 885 85
rect 885 15 905 85
rect 905 15 910 85
rect 880 10 910 15
rect 1130 85 1160 90
rect 1130 15 1135 85
rect 1135 15 1155 85
rect 1155 15 1160 85
rect 1130 10 1160 15
<< metal2 >>
rect 20 300 980 305
rect 20 220 25 300
rect 55 220 155 300
rect 185 220 430 300
rect 460 220 600 300
rect 630 220 650 300
rect 680 220 815 300
rect 845 220 945 300
rect 975 220 980 300
rect 20 215 980 220
rect -165 90 1165 95
rect -165 10 -160 90
rect -130 10 90 90
rect 120 10 430 90
rect 460 10 600 90
rect 630 10 650 90
rect 680 10 880 90
rect 910 10 1130 90
rect 1160 10 1165 90
rect -165 5 1165 10
<< end >>
