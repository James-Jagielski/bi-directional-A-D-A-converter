magic
tech sky130A
timestamp 1702662166
<< nwell >>
rect -90 595 0 715
rect -90 330 620 595
<< nmos >>
rect -20 150 -5 250
rect 45 150 60 250
rect 110 150 125 250
rect 175 150 190 250
rect 240 150 255 250
rect 385 150 400 250
rect -20 -165 -5 -65
rect 45 -165 60 -65
rect 110 -165 125 -65
rect 175 -165 190 -65
rect 240 -165 255 -65
rect 305 -165 320 -65
rect 370 -165 385 -65
<< pmos >>
rect -20 385 -5 485
rect 20 385 35 485
rect 85 385 100 485
rect 230 385 245 485
rect 295 385 310 485
rect 335 385 350 485
rect 480 385 495 485
<< ndiff >>
rect -70 235 -20 250
rect -70 165 -55 235
rect -35 165 -20 235
rect -70 150 -20 165
rect -5 235 45 250
rect -5 165 10 235
rect 30 165 45 235
rect -5 150 45 165
rect 60 235 110 250
rect 60 165 75 235
rect 95 165 110 235
rect 60 150 110 165
rect 125 235 175 250
rect 125 165 140 235
rect 160 165 175 235
rect 125 150 175 165
rect 190 235 240 250
rect 190 165 205 235
rect 225 165 240 235
rect 190 150 240 165
rect 255 235 305 250
rect 255 165 270 235
rect 290 165 305 235
rect 255 150 305 165
rect 335 235 385 250
rect 335 165 350 235
rect 370 165 385 235
rect 335 150 385 165
rect 400 235 450 250
rect 400 165 415 235
rect 435 165 450 235
rect 400 150 450 165
rect -70 -80 -20 -65
rect -70 -150 -55 -80
rect -35 -150 -20 -80
rect -70 -165 -20 -150
rect -5 -80 45 -65
rect -5 -150 10 -80
rect 30 -150 45 -80
rect -5 -165 45 -150
rect 60 -80 110 -65
rect 60 -150 75 -80
rect 95 -150 110 -80
rect 60 -165 110 -150
rect 125 -80 175 -65
rect 125 -150 140 -80
rect 160 -150 175 -80
rect 125 -165 175 -150
rect 190 -80 240 -65
rect 190 -150 205 -80
rect 225 -150 240 -80
rect 190 -165 240 -150
rect 255 -80 305 -65
rect 255 -150 270 -80
rect 290 -150 305 -80
rect 255 -165 305 -150
rect 320 -80 370 -65
rect 320 -150 335 -80
rect 355 -150 370 -80
rect 320 -165 370 -150
rect 385 -80 435 -65
rect 385 -150 400 -80
rect 420 -150 435 -80
rect 385 -165 435 -150
<< pdiff >>
rect -70 470 -20 485
rect -70 400 -55 470
rect -35 400 -20 470
rect -70 385 -20 400
rect -5 385 20 485
rect 35 470 85 485
rect 35 400 50 470
rect 70 400 85 470
rect 35 385 85 400
rect 100 470 150 485
rect 100 400 115 470
rect 135 400 150 470
rect 100 385 150 400
rect 180 470 230 485
rect 180 400 195 470
rect 215 400 230 470
rect 180 385 230 400
rect 245 470 295 485
rect 245 400 260 470
rect 280 400 295 470
rect 245 385 295 400
rect 310 385 335 485
rect 350 470 400 485
rect 350 400 365 470
rect 385 400 400 470
rect 350 385 400 400
rect 430 470 480 485
rect 430 400 445 470
rect 465 400 480 470
rect 430 385 480 400
rect 495 470 545 485
rect 495 400 510 470
rect 530 400 545 470
rect 495 385 545 400
<< ndiffc >>
rect -55 165 -35 235
rect 10 165 30 235
rect 75 165 95 235
rect 140 165 160 235
rect 205 165 225 235
rect 270 165 290 235
rect 350 165 370 235
rect 415 165 435 235
rect -55 -150 -35 -80
rect 10 -150 30 -80
rect 75 -150 95 -80
rect 140 -150 160 -80
rect 205 -150 225 -80
rect 270 -150 290 -80
rect 335 -150 355 -80
rect 400 -150 420 -80
<< pdiffc >>
rect -55 400 -35 470
rect 50 400 70 470
rect 115 400 135 470
rect 195 400 215 470
rect 260 400 280 470
rect 365 400 385 470
rect 445 400 465 470
rect 510 400 530 470
<< psubdiff >>
rect 475 -80 525 -65
rect 475 -150 490 -80
rect 510 -150 525 -80
rect 475 -165 525 -150
<< nsubdiff >>
rect -70 680 -20 695
rect -70 610 -55 680
rect -35 610 -20 680
rect -70 595 -20 610
<< psubdiffcont >>
rect 490 -150 510 -80
<< nsubdiffcont >>
rect -55 610 -35 680
<< poly >>
rect 100 530 140 540
rect 100 515 110 530
rect 20 510 110 515
rect 130 510 140 530
rect 20 500 140 510
rect 190 530 230 540
rect 190 510 200 530
rect 220 515 230 530
rect 335 525 640 540
rect 220 510 310 515
rect 190 500 310 510
rect -20 485 -5 500
rect 20 485 35 500
rect 85 485 100 500
rect 230 485 245 500
rect 295 485 310 500
rect 335 485 350 525
rect 480 485 495 500
rect -20 345 -5 385
rect 20 370 35 385
rect 85 370 100 385
rect 230 370 245 385
rect 295 370 310 385
rect 335 345 350 385
rect -135 330 350 345
rect 45 290 255 305
rect 45 280 60 290
rect -135 265 60 280
rect -20 250 -5 265
rect 45 250 60 265
rect 110 250 125 265
rect 175 250 190 265
rect 240 250 255 290
rect 385 250 400 265
rect -20 135 -5 150
rect 45 135 60 150
rect 110 110 125 150
rect -135 95 125 110
rect 175 70 190 150
rect 240 135 255 150
rect 385 135 400 150
rect 480 135 495 385
rect 385 125 425 135
rect 385 105 395 125
rect 415 105 425 125
rect 385 95 425 105
rect 455 125 495 135
rect 455 105 465 125
rect 485 105 495 125
rect 455 95 495 105
rect 580 285 645 305
rect 580 70 600 285
rect 175 55 600 70
rect 630 30 670 40
rect 45 20 640 30
rect 45 15 455 20
rect -135 -50 -5 -35
rect -20 -65 -5 -50
rect 45 -65 60 15
rect 175 -20 215 -10
rect 175 -40 185 -20
rect 205 -40 215 -20
rect 175 -50 215 -40
rect 300 -20 340 -10
rect 300 -40 310 -20
rect 330 -40 340 -20
rect 300 -50 340 -40
rect 110 -65 125 -50
rect 175 -65 190 -50
rect 240 -65 255 -50
rect 305 -65 320 -50
rect 370 -65 385 15
rect 445 0 455 15
rect 475 15 640 20
rect 475 0 485 15
rect 630 10 640 15
rect 660 10 670 30
rect 630 0 670 10
rect 445 -10 485 0
rect -20 -180 -5 -165
rect 45 -180 60 -165
rect 110 -245 125 -165
rect 175 -180 190 -165
rect 150 -190 190 -180
rect 150 -210 160 -190
rect 180 -210 190 -190
rect 150 -220 190 -210
rect 240 -180 255 -165
rect 305 -180 320 -165
rect 370 -180 385 -165
rect 240 -190 280 -180
rect 240 -210 250 -190
rect 270 -210 280 -190
rect 240 -220 280 -210
rect 110 -260 645 -245
<< polycont >>
rect 110 510 130 530
rect 200 510 220 530
rect 395 105 415 125
rect 465 105 485 125
rect 185 -40 205 -20
rect 310 -40 330 -20
rect 455 0 475 20
rect 640 10 660 30
rect 160 -210 180 -190
rect 250 -210 270 -190
<< locali >>
rect -65 680 -25 690
rect -65 610 -55 680
rect -35 610 -25 680
rect -65 600 -25 610
rect 575 590 615 595
rect 575 580 585 590
rect -45 570 585 580
rect 605 580 615 590
rect 605 570 640 580
rect -45 560 640 570
rect -45 480 -25 560
rect 100 530 140 540
rect 100 510 110 530
rect 130 510 140 530
rect 100 500 140 510
rect 190 530 230 540
rect 190 510 200 530
rect 220 510 230 530
rect 190 500 230 510
rect 375 500 640 520
rect 105 480 125 500
rect 205 480 225 500
rect 375 480 395 500
rect -65 470 -25 480
rect -65 400 -55 470
rect -35 400 -25 470
rect -65 390 -25 400
rect 40 470 80 480
rect 40 400 50 470
rect 70 400 80 470
rect 40 390 80 400
rect 105 470 145 480
rect 105 400 115 470
rect 135 400 145 470
rect 105 390 145 400
rect 125 360 145 390
rect 85 340 145 360
rect 185 470 225 480
rect 185 400 195 470
rect 215 400 225 470
rect 185 390 225 400
rect 250 470 290 480
rect 250 400 260 470
rect 280 400 290 470
rect 250 390 290 400
rect 355 470 395 480
rect 355 400 365 470
rect 385 400 395 470
rect 355 390 395 400
rect 435 470 475 480
rect 435 400 445 470
rect 465 400 475 470
rect 435 390 475 400
rect 500 470 540 480
rect 500 400 510 470
rect 530 400 540 470
rect 500 390 540 400
rect 185 360 205 390
rect 375 375 395 390
rect 185 340 215 360
rect 375 355 425 375
rect 85 245 105 340
rect 195 245 215 340
rect 405 245 425 355
rect -65 235 -25 245
rect -65 165 -55 235
rect -35 165 -25 235
rect -65 155 -25 165
rect 0 235 40 245
rect 0 165 10 235
rect 30 165 40 235
rect 0 155 40 165
rect 65 235 105 245
rect 65 165 75 235
rect 95 165 105 235
rect 65 155 105 165
rect 130 235 170 245
rect 130 165 140 235
rect 160 165 170 235
rect 130 155 170 165
rect 195 235 235 245
rect 195 165 205 235
rect 225 165 235 235
rect 195 155 235 165
rect 260 235 300 245
rect 260 165 270 235
rect 290 165 300 235
rect 260 155 300 165
rect 340 235 380 245
rect 340 165 350 235
rect 370 165 380 235
rect 340 155 380 165
rect 405 235 445 245
rect 405 165 415 235
rect 435 165 445 235
rect 405 155 445 165
rect -45 135 -25 155
rect 130 135 150 155
rect -45 115 150 135
rect 340 40 360 155
rect 385 125 425 135
rect 385 105 395 125
rect 415 105 425 125
rect 385 95 425 105
rect 455 125 495 135
rect 455 105 465 125
rect 485 105 495 125
rect 455 95 495 105
rect 130 20 360 40
rect 130 -70 150 20
rect 175 -20 215 -10
rect 175 -40 185 -20
rect 205 -30 215 -20
rect 300 -20 340 -10
rect 205 -40 280 -30
rect 175 -50 280 -40
rect 300 -40 310 -20
rect 330 -30 340 -20
rect 390 -30 410 95
rect 465 30 485 95
rect 445 20 485 30
rect 445 0 455 20
rect 475 0 485 20
rect 445 -10 485 0
rect 520 -30 540 390
rect 330 -40 540 -30
rect 300 -50 540 -40
rect 580 465 620 475
rect 580 445 590 465
rect 610 445 620 465
rect 580 435 620 445
rect 260 -70 280 -50
rect 390 -70 410 -50
rect -65 -80 -25 -70
rect -65 -150 -55 -80
rect -35 -150 -25 -80
rect -65 -170 -25 -150
rect 0 -80 40 -70
rect 0 -150 10 -80
rect 30 -150 40 -80
rect 0 -160 40 -150
rect -65 -190 -55 -170
rect -35 -190 -25 -170
rect -65 -200 -25 -190
rect -45 -260 -25 -200
rect 20 -220 40 -160
rect 65 -80 105 -70
rect 65 -150 75 -80
rect 95 -150 105 -80
rect 65 -170 105 -150
rect 130 -80 170 -70
rect 130 -150 140 -80
rect 160 -150 170 -80
rect 130 -160 170 -150
rect 195 -80 235 -70
rect 195 -150 205 -80
rect 225 -150 235 -80
rect 195 -160 235 -150
rect 260 -80 300 -70
rect 260 -150 270 -80
rect 290 -150 300 -80
rect 260 -160 300 -150
rect 325 -80 365 -70
rect 325 -150 335 -80
rect 355 -150 365 -80
rect 325 -160 365 -150
rect 390 -80 430 -70
rect 390 -150 400 -80
rect 420 -150 430 -80
rect 390 -160 430 -150
rect 480 -80 520 -70
rect 480 -150 490 -80
rect 510 -150 520 -80
rect 480 -160 520 -150
rect 65 -190 75 -170
rect 95 -190 105 -170
rect 345 -180 365 -160
rect 580 -180 600 435
rect 630 30 670 40
rect 630 10 640 30
rect 660 10 670 30
rect 630 0 670 10
rect 65 -200 105 -190
rect 150 -190 190 -180
rect 150 -210 160 -190
rect 180 -210 190 -190
rect 150 -220 190 -210
rect 240 -190 280 -180
rect 240 -210 250 -190
rect 270 -210 280 -190
rect 345 -200 600 -180
rect 240 -220 280 -210
rect 20 -240 170 -220
rect 240 -260 260 -220
rect -45 -280 260 -260
<< viali >>
rect -55 610 -35 680
rect 585 570 605 590
rect 50 400 70 470
rect 260 400 280 470
rect 445 400 465 470
rect 10 165 30 235
rect 270 165 290 235
rect 590 445 610 465
rect -55 -190 -35 -170
rect 205 -150 225 -80
rect 490 -150 510 -80
rect 75 -190 95 -170
<< metal1 >>
rect -65 685 -25 690
rect -65 605 -60 685
rect -30 605 -25 685
rect -65 600 -25 605
rect 575 590 615 595
rect 575 570 585 590
rect 605 570 615 590
rect 575 560 615 570
rect 40 475 80 480
rect 40 395 45 475
rect 75 395 80 475
rect 40 390 80 395
rect 250 475 290 480
rect 250 395 255 475
rect 285 395 290 475
rect 250 390 290 395
rect 435 475 475 480
rect 435 395 440 475
rect 470 395 475 475
rect 580 475 600 560
rect 580 465 620 475
rect 580 445 590 465
rect 610 445 620 465
rect 580 435 620 445
rect 435 390 475 395
rect 0 240 40 250
rect 0 160 5 240
rect 35 160 40 240
rect 0 150 40 160
rect 255 240 305 250
rect 255 160 265 240
rect 295 160 305 240
rect 255 150 305 160
rect 190 -75 240 -65
rect 190 -155 200 -75
rect 230 -155 240 -75
rect -65 -170 105 -160
rect 190 -165 240 -155
rect 480 -75 520 -70
rect 480 -155 485 -75
rect 515 -155 520 -75
rect 480 -160 520 -155
rect -65 -190 -55 -170
rect -35 -190 75 -170
rect 95 -190 105 -170
rect -65 -200 105 -190
<< via1 >>
rect -60 680 -30 685
rect -60 610 -55 680
rect -55 610 -35 680
rect -35 610 -30 680
rect -60 605 -30 610
rect 45 470 75 475
rect 45 400 50 470
rect 50 400 70 470
rect 70 400 75 470
rect 45 395 75 400
rect 255 470 285 475
rect 255 400 260 470
rect 260 400 280 470
rect 280 400 285 470
rect 255 395 285 400
rect 440 470 470 475
rect 440 400 445 470
rect 445 400 465 470
rect 465 400 470 470
rect 440 395 470 400
rect 5 235 35 240
rect 5 165 10 235
rect 10 165 30 235
rect 30 165 35 235
rect 5 160 35 165
rect 265 235 295 240
rect 265 165 270 235
rect 270 165 290 235
rect 290 165 295 235
rect 265 160 295 165
rect 200 -80 230 -75
rect 200 -150 205 -80
rect 205 -150 225 -80
rect 225 -150 230 -80
rect 200 -155 230 -150
rect 485 -80 515 -75
rect 485 -150 490 -80
rect 490 -150 510 -80
rect 510 -150 515 -80
rect 485 -155 515 -150
<< metal2 >>
rect -70 685 -20 695
rect -70 605 -60 685
rect -30 605 -20 685
rect -70 595 -20 605
rect -70 480 550 595
rect -70 475 545 480
rect -70 395 45 475
rect 75 395 255 475
rect 285 395 440 475
rect 470 395 545 475
rect -70 390 545 395
rect -115 240 620 255
rect -115 160 5 240
rect 35 160 265 240
rect 295 160 620 240
rect -115 70 620 160
rect -135 55 620 70
rect -115 -75 620 55
rect -115 -155 200 -75
rect 230 -155 485 -75
rect 515 -155 620 -75
rect -115 -160 620 -155
<< labels >>
rlabel poly -135 100 -135 100 7 AIn
port 1 w
rlabel poly -135 -45 -135 -45 7 RST
port 2 w
rlabel poly 645 -255 645 -255 3 ENAD
port 3 e
rlabel locali 640 570 640 570 3 CompOut
port 6 e
rlabel poly -135 270 -135 270 7 Vb
port 7 w
<< end >>
