magic
tech sky130A
timestamp 1702693377
<< nwell >>
rect 170 2170 345 2310
<< nmos >>
rect 240 2035 255 2135
<< pmos >>
rect 240 2190 255 2290
<< ndiff >>
rect 190 2120 240 2135
rect 190 2050 205 2120
rect 225 2050 240 2120
rect 190 2035 240 2050
rect 255 2120 305 2135
rect 255 2050 270 2120
rect 290 2050 305 2120
rect 255 2035 305 2050
<< pdiff >>
rect 190 2275 240 2290
rect 190 2205 205 2275
rect 225 2205 240 2275
rect 190 2190 240 2205
rect 255 2275 305 2290
rect 255 2205 270 2275
rect 290 2205 305 2275
rect 255 2190 305 2205
<< ndiffc >>
rect 205 2050 225 2120
rect 270 2050 290 2120
<< pdiffc >>
rect 205 2205 225 2275
rect 270 2205 290 2275
<< poly >>
rect 2455 3370 2495 3380
rect 2455 3350 2465 3370
rect 2485 3350 2495 3370
rect 2455 3340 2495 3350
rect 2635 3340 2665 3370
rect 1050 3110 1090 3120
rect 1050 3095 1060 3110
rect 1005 3090 1060 3095
rect 1080 3090 1090 3110
rect 140 3070 180 3080
rect 1005 3075 1090 3090
rect 140 3050 150 3070
rect 170 3055 270 3070
rect 170 3050 180 3055
rect 140 3045 180 3050
rect 155 3040 180 3045
rect 2340 2935 2380 2945
rect 2340 2915 2350 2935
rect 2370 2915 2380 2935
rect 45 2900 85 2910
rect 2340 2905 2380 2915
rect 45 2880 55 2900
rect 75 2885 270 2900
rect 75 2880 85 2885
rect 45 2870 85 2880
rect 1865 2865 1905 2875
rect 1865 2845 1875 2865
rect 1895 2845 1905 2865
rect 1865 2835 1905 2845
rect 2155 2870 2195 2880
rect 2155 2850 2165 2870
rect 2185 2850 2195 2870
rect 2155 2840 2195 2850
rect 1410 2825 1450 2835
rect 1410 2805 1420 2825
rect 1440 2810 1450 2825
rect 2465 2810 2485 3340
rect 1440 2805 2485 2810
rect 1410 2795 2485 2805
rect 50 2760 90 2770
rect 50 2740 60 2760
rect 80 2755 90 2760
rect 80 2740 250 2755
rect 50 2730 90 2740
rect -95 2550 -55 2560
rect -95 2530 -85 2550
rect -65 2545 -55 2550
rect -65 2530 665 2545
rect -95 2520 -55 2530
rect 715 2480 755 2490
rect 715 2460 725 2480
rect 745 2460 755 2480
rect 715 2450 755 2460
rect 280 2335 320 2345
rect 280 2315 290 2335
rect 310 2320 320 2335
rect 310 2315 405 2320
rect 280 2305 405 2315
rect 240 2290 255 2305
rect 2342 2266 2382 2274
rect 2342 2247 2354 2266
rect 2373 2253 2382 2266
rect 2555 2259 2598 2270
rect 2555 2253 2567 2259
rect 2373 2247 2567 2253
rect 2342 2241 2567 2247
rect 2586 2241 2598 2259
rect 2342 2236 2598 2241
rect 2342 2235 2382 2236
rect 2555 2226 2598 2236
rect 240 2135 255 2190
rect -110 2005 -70 2015
rect -110 1985 -100 2005
rect -80 2000 -70 2005
rect 240 2000 255 2035
rect -80 1985 255 2000
rect -110 1980 255 1985
rect -110 1975 -70 1980
rect 240 1665 255 1980
rect 300 1930 405 1950
rect 2575 1945 2615 1955
rect 300 1730 320 1930
rect 2265 1925 2585 1945
rect 2605 1925 2615 1945
rect 2575 1915 2615 1925
rect 1379 1815 1416 1824
rect 1379 1796 1387 1815
rect 1405 1796 1416 1815
rect 1379 1790 1416 1796
rect 1295 1763 1310 1772
rect 1382 1763 1399 1790
rect 1295 1744 1399 1763
rect 295 1725 335 1730
rect 295 1700 300 1725
rect 325 1700 335 1725
rect 295 1690 335 1700
rect 240 1650 420 1665
<< polycont >>
rect 2465 3350 2485 3370
rect 1060 3090 1080 3110
rect 150 3050 170 3070
rect 2350 2915 2370 2935
rect 55 2880 75 2900
rect 1875 2845 1895 2865
rect 2165 2850 2185 2870
rect 1420 2805 1440 2825
rect 60 2740 80 2760
rect -85 2530 -65 2550
rect 725 2460 745 2480
rect 290 2315 310 2335
rect 2354 2247 2373 2266
rect 2567 2241 2586 2259
rect -100 1985 -80 2005
rect 2585 1925 2605 1945
rect 1387 1796 1405 1815
rect 300 1700 325 1725
<< locali >>
rect 1610 3463 1662 3474
rect 1610 3437 1624 3463
rect 1650 3437 1662 3463
rect 1610 3425 1662 3437
rect 1630 3344 1650 3425
rect 2005 3375 2045 3385
rect 2005 3355 2015 3375
rect 2035 3355 2045 3375
rect 2005 3345 2045 3355
rect 2255 3370 2295 3380
rect 2255 3350 2265 3370
rect 2285 3350 2295 3370
rect 2010 3265 2030 3345
rect 2255 3340 2295 3350
rect 2455 3370 2495 3380
rect 2455 3350 2465 3370
rect 2485 3350 2495 3370
rect 2455 3340 2495 3350
rect 2635 3340 2665 3370
rect 2260 3255 2280 3340
rect 1050 3110 1090 3120
rect 2310 3115 2325 3140
rect 1050 3090 1060 3110
rect 1080 3090 1090 3110
rect 1050 3080 1090 3090
rect 140 3070 180 3080
rect 140 3050 150 3070
rect 170 3050 180 3070
rect 140 3045 180 3050
rect 1165 2935 1185 2995
rect 1150 2925 1190 2935
rect 45 2900 85 2910
rect 45 2880 55 2900
rect 75 2880 85 2900
rect 1150 2905 1160 2925
rect 1180 2905 1190 2925
rect 1150 2895 1190 2905
rect 45 2870 85 2880
rect 1790 2865 1810 2980
rect 1865 2865 1905 2875
rect 1790 2845 1875 2865
rect 1895 2845 1905 2865
rect 1865 2835 1905 2845
rect 1410 2825 1450 2835
rect 1410 2805 1420 2825
rect 1440 2805 1450 2825
rect 1410 2795 1450 2805
rect 2010 2820 2030 2980
rect 2155 2870 2195 2880
rect 2155 2850 2165 2870
rect 2185 2850 2195 2870
rect 2155 2840 2195 2850
rect 2295 2875 2315 2985
rect 2340 2935 2380 2945
rect 2340 2915 2350 2935
rect 2370 2915 2380 2935
rect 2340 2905 2380 2915
rect 2295 2845 2425 2875
rect 2010 2800 2320 2820
rect 50 2760 90 2770
rect 50 2740 60 2760
rect 80 2740 90 2760
rect 50 2730 90 2740
rect -95 2550 -55 2560
rect -95 2530 -85 2550
rect -65 2530 -55 2550
rect -95 2520 -55 2530
rect 715 2480 755 2490
rect 715 2460 725 2480
rect 745 2460 755 2480
rect 715 2450 755 2460
rect -100 2400 -60 2410
rect 200 2405 245 2415
rect 1415 2405 1435 2795
rect 200 2400 210 2405
rect -100 2380 -90 2400
rect -70 2380 210 2400
rect 235 2380 245 2405
rect -100 2375 245 2380
rect -100 2370 -60 2375
rect 200 2370 245 2375
rect 280 2335 320 2345
rect 280 2315 290 2335
rect 310 2315 320 2335
rect 2290 2325 2320 2800
rect 280 2305 320 2315
rect 2125 2305 2320 2325
rect 280 2285 300 2305
rect 200 2275 235 2285
rect 200 2205 205 2275
rect 225 2205 235 2275
rect 200 2195 235 2205
rect 260 2275 300 2285
rect 260 2205 270 2275
rect 290 2205 300 2275
rect 2342 2266 2382 2274
rect 2342 2249 2354 2266
rect 2337 2247 2354 2249
rect 2373 2247 2382 2266
rect 2337 2235 2382 2247
rect 2337 2214 2359 2235
rect -111 2148 -71 2159
rect -111 2127 -102 2148
rect -81 2138 -71 2148
rect -81 2127 10 2138
rect -111 2119 10 2127
rect -111 2117 -71 2119
rect -110 2005 -70 2015
rect -110 1985 -100 2005
rect -80 1985 -70 2005
rect -110 1975 -70 1985
rect -12 2002 10 2119
rect 200 2120 235 2130
rect 200 2050 205 2120
rect 225 2050 235 2120
rect 200 2040 235 2050
rect 260 2120 300 2205
rect 260 2050 270 2120
rect 290 2050 300 2120
rect 260 2040 300 2050
rect -12 1980 340 2002
rect -10 1979 340 1980
rect -115 1895 -70 1905
rect -115 1875 -105 1895
rect -85 1875 -70 1895
rect -115 1865 -70 1875
rect 320 1865 340 1895
rect -100 1730 -70 1865
rect 1379 1815 1416 1824
rect 1379 1795 1385 1815
rect 1406 1795 1416 1815
rect 1379 1790 1416 1795
rect -100 1725 335 1730
rect -100 1705 300 1725
rect 295 1700 300 1705
rect 325 1700 335 1725
rect 2400 1710 2425 2845
rect 2555 2259 2598 2270
rect 2555 2241 2567 2259
rect 2586 2241 2598 2259
rect 2555 2226 2598 2241
rect 2575 1945 2615 1955
rect 2575 1925 2585 1945
rect 2605 1925 2615 1945
rect 2575 1915 2615 1925
rect 295 1690 335 1700
rect 2105 1690 2425 1710
rect 155 1600 175 1605
rect 2350 810 2390 820
rect 2350 790 2360 810
rect 2380 790 2390 810
rect 2350 780 2390 790
<< viali >>
rect 1624 3437 1650 3463
rect 2015 3355 2035 3375
rect 2265 3350 2285 3370
rect 2465 3350 2485 3370
rect 1060 3090 1080 3110
rect 150 3050 170 3070
rect 1470 2975 1490 3045
rect 55 2880 75 2900
rect 1160 2905 1180 2925
rect 1320 2915 1340 2935
rect 1875 2845 1895 2865
rect 1420 2805 1440 2825
rect 2165 2850 2185 2870
rect 2350 2915 2370 2935
rect 60 2740 80 2760
rect 550 2750 570 2770
rect 615 2580 635 2600
rect -85 2530 -65 2550
rect 725 2460 745 2480
rect -90 2380 -70 2400
rect 210 2380 235 2405
rect 1690 2315 1710 2335
rect 205 2205 225 2275
rect 1605 2205 1625 2275
rect -102 2127 -81 2148
rect -100 1985 -80 2005
rect 205 2050 225 2120
rect -105 1875 -85 1895
rect 1385 1796 1387 1815
rect 1387 1796 1405 1815
rect 1405 1796 1406 1815
rect 1385 1795 1406 1796
rect 1060 1700 1080 1720
rect 2567 2241 2586 2259
rect 2585 1925 2605 1945
rect 300 1595 320 1615
rect 2360 1600 2380 1620
rect 2360 790 2380 810
<< metal1 >>
rect -11 3644 796 3669
rect -11 2910 14 3644
rect 769 3460 794 3644
rect 1610 3463 1662 3474
rect 1610 3460 1624 3463
rect 535 3455 575 3460
rect 535 3425 540 3455
rect 570 3425 575 3455
rect 535 3420 575 3425
rect 620 3455 660 3460
rect 620 3425 625 3455
rect 655 3440 660 3455
rect 655 3425 715 3440
rect 769 3437 1624 3460
rect 1650 3437 1662 3463
rect 769 3436 794 3437
rect 1610 3425 1662 3437
rect 620 3420 715 3425
rect 140 3070 180 3080
rect 140 3050 150 3070
rect 170 3050 180 3070
rect 140 3040 180 3050
rect -11 2900 85 2910
rect -11 2880 55 2900
rect 75 2880 85 2900
rect -11 2878 14 2880
rect 45 2870 85 2880
rect 50 2765 90 2770
rect -1000 2760 90 2765
rect -1000 2740 60 2760
rect 80 2740 90 2760
rect 50 2730 90 2740
rect -1000 2550 -55 2560
rect -1000 2535 -85 2550
rect -95 2530 -85 2535
rect -65 2530 -55 2550
rect -95 2520 -55 2530
rect -100 2405 -60 2410
rect -100 2375 -95 2405
rect -65 2375 -60 2405
rect -100 2370 -60 2375
rect -1003 2148 -71 2159
rect -1003 2132 -102 2148
rect -111 2127 -102 2132
rect -81 2127 -71 2148
rect -111 2117 -71 2127
rect -110 2005 -70 2015
rect -110 2000 -100 2005
rect -1000 1985 -100 2000
rect -80 1985 -70 2005
rect -1000 1975 -70 1985
rect -115 1900 -75 1905
rect -115 1870 -110 1900
rect -80 1870 -75 1900
rect -115 1865 -75 1870
rect -1000 1689 -899 1690
rect 86 1689 123 1698
rect -1000 1667 123 1689
rect -1000 1666 -899 1667
rect 86 1658 123 1667
rect 155 1625 180 3040
rect 540 2780 560 3420
rect 625 3180 645 3275
rect 625 2940 645 3035
rect 695 2905 715 3420
rect 2005 3380 2045 3385
rect 2005 3350 2010 3380
rect 2040 3350 2045 3380
rect 2005 3345 2045 3350
rect 2255 3375 2295 3380
rect 2255 3345 2260 3375
rect 2290 3345 2295 3375
rect 2255 3340 2295 3345
rect 2455 3375 2495 3380
rect 2455 3345 2460 3375
rect 2490 3345 2495 3375
rect 2455 3340 2495 3345
rect 2630 3370 2670 3375
rect 2630 3340 2635 3370
rect 2665 3340 2670 3370
rect 2630 3335 2670 3340
rect 1610 3125 1635 3130
rect 1050 3115 2610 3125
rect 1050 3110 2575 3115
rect 1050 3090 1060 3110
rect 1080 3090 2575 3110
rect 1050 3085 2575 3090
rect 2605 3085 2610 3115
rect 1050 3080 2610 3085
rect 1460 3045 1500 3055
rect 1460 2975 1470 3045
rect 1490 2975 1500 3045
rect 1460 2965 1500 2975
rect 1310 2935 1350 2945
rect 625 2885 715 2905
rect 1150 2930 1190 2935
rect 1150 2900 1155 2930
rect 1185 2900 1190 2930
rect 1310 2915 1320 2935
rect 1340 2930 1350 2935
rect 1340 2915 1385 2930
rect 1310 2910 1385 2915
rect 1310 2905 1350 2910
rect 1150 2895 1190 2900
rect 540 2770 580 2780
rect 540 2750 550 2770
rect 570 2750 580 2770
rect 540 2740 580 2750
rect 625 2610 645 2885
rect 605 2600 645 2610
rect 605 2580 615 2600
rect 635 2580 645 2600
rect 605 2570 645 2580
rect 1365 2660 1385 2910
rect 1470 2835 1490 2965
rect 1410 2825 1490 2835
rect 1410 2805 1420 2825
rect 1440 2820 1490 2825
rect 1440 2815 1485 2820
rect 1440 2805 1450 2815
rect 1410 2795 1450 2805
rect 1610 2795 1635 3080
rect 2635 2945 2665 3335
rect 2340 2935 2380 2945
rect 2340 2915 2350 2935
rect 2370 2915 2380 2935
rect 1865 2865 1905 2875
rect 1865 2845 1875 2865
rect 1895 2845 1905 2865
rect 1865 2835 1905 2845
rect 2155 2870 2195 2880
rect 2155 2850 2165 2870
rect 2185 2850 2195 2870
rect 2155 2840 2195 2850
rect 1605 2790 1645 2795
rect 1605 2760 1610 2790
rect 1640 2760 1645 2790
rect 1605 2755 1645 2760
rect 1405 2730 1450 2735
rect 1865 2730 1885 2835
rect 2170 2765 2195 2840
rect 1405 2700 1415 2730
rect 1445 2710 1885 2730
rect 2155 2760 2195 2765
rect 2155 2730 2160 2760
rect 2190 2730 2195 2760
rect 2155 2725 2195 2730
rect 1445 2700 1450 2710
rect 1405 2695 1450 2700
rect 2155 2660 2195 2665
rect 1365 2640 2160 2660
rect 715 2485 755 2490
rect 1365 2485 1385 2640
rect 1410 2585 1870 2595
rect 1410 2555 1415 2585
rect 1445 2575 1870 2585
rect 1445 2555 1450 2575
rect 1410 2550 1450 2555
rect 1605 2515 1645 2520
rect 715 2455 720 2485
rect 750 2455 755 2485
rect 715 2450 755 2455
rect 825 2460 1385 2485
rect 1410 2510 1450 2515
rect 1410 2480 1415 2510
rect 1445 2480 1450 2510
rect 1605 2485 1610 2515
rect 1640 2485 1645 2515
rect 1605 2480 1645 2485
rect 1410 2475 1450 2480
rect 200 2410 245 2415
rect 200 2375 205 2410
rect 240 2375 245 2410
rect 200 2370 245 2375
rect 195 2280 235 2285
rect 195 2200 200 2280
rect 230 2200 235 2280
rect 195 2195 235 2200
rect 195 2125 235 2130
rect 195 2045 200 2125
rect 230 2045 235 2125
rect 195 2040 235 2045
rect 290 2120 510 2160
rect 290 1625 330 2120
rect 725 2100 750 2450
rect 825 2130 845 2460
rect 880 2405 920 2410
rect 880 2375 885 2405
rect 915 2390 1305 2405
rect 915 2375 920 2390
rect 880 2370 920 2375
rect 1290 2285 1305 2390
rect 1381 1824 1401 1825
rect 1379 1815 1416 1824
rect 1379 1795 1385 1815
rect 1406 1795 1416 1815
rect 1379 1790 1416 1795
rect 1381 1769 1401 1790
rect 1362 1766 1406 1769
rect 1050 1720 1090 1730
rect 1362 1729 1366 1766
rect 1401 1729 1406 1766
rect 1362 1726 1406 1729
rect 1050 1700 1060 1720
rect 1080 1710 1090 1720
rect 1430 1710 1445 2475
rect 1610 2285 1635 2480
rect 1680 2340 1720 2345
rect 1680 2310 1685 2340
rect 1715 2310 1720 2340
rect 1680 2305 1720 2310
rect 1590 2275 1635 2285
rect 1590 2205 1605 2275
rect 1625 2205 1635 2275
rect 1590 2195 1635 2205
rect 1850 2110 1870 2575
rect 1910 2100 1935 2640
rect 2155 2630 2160 2640
rect 2190 2630 2195 2660
rect 2155 2625 2195 2630
rect 2340 2345 2380 2915
rect 2430 2940 2665 2945
rect 2430 2910 2435 2940
rect 2465 2920 2665 2940
rect 2465 2910 2470 2920
rect 2430 2905 2470 2910
rect 2440 2760 2480 2765
rect 2440 2755 2445 2760
rect 2430 2735 2445 2755
rect 2440 2730 2445 2735
rect 2475 2755 2480 2760
rect 2475 2735 3725 2755
rect 2475 2730 2480 2735
rect 2440 2725 2480 2730
rect 2440 2660 2480 2665
rect 2440 2630 2445 2660
rect 2475 2655 2480 2660
rect 2475 2635 3725 2655
rect 2475 2630 2480 2635
rect 2440 2625 2480 2630
rect 2230 2340 2445 2345
rect 2230 2310 2235 2340
rect 2265 2310 2445 2340
rect 2230 2305 2445 2310
rect 2165 2120 2390 2160
rect 1080 1700 1445 1710
rect 1050 1690 1445 1700
rect 155 1615 330 1625
rect 155 1595 300 1615
rect 320 1595 330 1615
rect 155 1585 330 1595
rect 2350 1620 2390 2120
rect 2405 1680 2445 2305
rect 2558 2259 2598 2269
rect 2558 2241 2567 2259
rect 2586 2244 2598 2259
rect 2586 2241 3746 2244
rect 2558 2225 3746 2241
rect 2575 1950 2615 1955
rect 2575 1920 2580 1950
rect 2610 1920 2615 1950
rect 2575 1915 2615 1920
rect 2405 1640 2645 1680
rect 2350 1600 2360 1620
rect 2380 1600 2390 1620
rect 2350 1590 2390 1600
rect 2605 820 2645 1640
rect 2350 810 2645 820
rect 2350 790 2360 810
rect 2380 790 2645 810
rect 2350 780 2645 790
<< via1 >>
rect 540 3425 570 3455
rect 625 3425 655 3455
rect -95 2400 -65 2405
rect -95 2380 -90 2400
rect -90 2380 -70 2400
rect -70 2380 -65 2400
rect -95 2375 -65 2380
rect -110 1895 -80 1900
rect -110 1875 -105 1895
rect -105 1875 -85 1895
rect -85 1875 -80 1895
rect -110 1870 -80 1875
rect 2010 3375 2040 3380
rect 2010 3355 2015 3375
rect 2015 3355 2035 3375
rect 2035 3355 2040 3375
rect 2010 3350 2040 3355
rect 2260 3370 2290 3375
rect 2260 3350 2265 3370
rect 2265 3350 2285 3370
rect 2285 3350 2290 3370
rect 2260 3345 2290 3350
rect 2460 3370 2490 3375
rect 2460 3350 2465 3370
rect 2465 3350 2485 3370
rect 2485 3350 2490 3370
rect 2460 3345 2490 3350
rect 2635 3340 2665 3370
rect 2575 3085 2605 3115
rect 1155 2925 1185 2930
rect 1155 2905 1160 2925
rect 1160 2905 1180 2925
rect 1180 2905 1185 2925
rect 1155 2900 1185 2905
rect 1610 2760 1640 2790
rect 1415 2700 1445 2730
rect 2160 2730 2190 2760
rect 1415 2555 1445 2585
rect 720 2480 750 2485
rect 720 2460 725 2480
rect 725 2460 745 2480
rect 745 2460 750 2480
rect 720 2455 750 2460
rect 1415 2480 1445 2510
rect 1610 2485 1640 2515
rect 205 2405 240 2410
rect 205 2380 210 2405
rect 210 2380 235 2405
rect 235 2380 240 2405
rect 205 2375 240 2380
rect 200 2275 230 2280
rect 200 2205 205 2275
rect 205 2205 225 2275
rect 225 2205 230 2275
rect 200 2200 230 2205
rect 200 2120 230 2125
rect 200 2050 205 2120
rect 205 2050 225 2120
rect 225 2050 230 2120
rect 200 2045 230 2050
rect 885 2375 915 2405
rect 1366 1729 1401 1766
rect 1685 2335 1715 2340
rect 1685 2315 1690 2335
rect 1690 2315 1710 2335
rect 1710 2315 1715 2335
rect 1685 2310 1715 2315
rect 2160 2630 2190 2660
rect 2435 2910 2465 2940
rect 2445 2730 2475 2760
rect 2445 2630 2475 2660
rect 2235 2310 2265 2340
rect 2580 1945 2610 1950
rect 2580 1925 2585 1945
rect 2585 1925 2605 1945
rect 2605 1925 2610 1945
rect 2580 1920 2610 1925
<< metal2 >>
rect -885 5210 -880 5240
rect -850 5210 -845 5240
rect -885 4425 -845 5210
rect -110 5210 -105 5240
rect -75 5210 -70 5240
rect -110 4660 -70 5210
rect 665 5210 670 5240
rect 700 5210 705 5240
rect -110 4630 650 4660
rect -885 4405 565 4425
rect -1015 3385 365 3505
rect 545 3460 565 4405
rect 630 3460 650 4630
rect 665 4425 705 5210
rect 1440 5210 1445 5240
rect 1475 5210 1480 5240
rect 1440 4470 1480 5210
rect 2215 5210 2220 5240
rect 2250 5210 2255 5240
rect 2215 4485 2255 5210
rect 2990 5210 2995 5240
rect 3025 5210 3030 5240
rect 1440 4450 2170 4470
rect 2215 4455 2480 4485
rect 665 4410 2030 4425
rect 535 3455 575 3460
rect 535 3425 540 3455
rect 570 3425 575 3455
rect 535 3420 575 3425
rect 620 3455 660 3460
rect 620 3425 625 3455
rect 655 3425 660 3455
rect 620 3420 660 3425
rect 2010 3385 2030 4410
rect 2145 4420 2170 4450
rect 2145 4405 2280 4420
rect 2005 3380 2045 3385
rect 2260 3380 2280 4405
rect 2460 3380 2480 4455
rect 2990 4425 3030 5210
rect 2635 4400 3030 4425
rect 2005 3350 2010 3380
rect 2040 3350 2045 3380
rect 2005 3345 2045 3350
rect 2255 3375 2295 3380
rect 2255 3345 2260 3375
rect 2290 3345 2295 3375
rect 2255 3340 2295 3345
rect 2455 3375 2495 3380
rect 2635 3375 2655 4400
rect 2455 3345 2460 3375
rect 2490 3345 2495 3375
rect 2455 3340 2495 3345
rect 2630 3370 2670 3375
rect 2630 3340 2635 3370
rect 2665 3340 2670 3370
rect 2630 3335 2670 3340
rect 2185 3175 2550 3230
rect 2430 2940 2470 2945
rect 1150 2930 1190 2935
rect 1150 2900 1155 2930
rect 1185 2900 1190 2930
rect 1150 2895 1190 2900
rect 1165 2885 1190 2895
rect 2430 2910 2435 2940
rect 2465 2910 2470 2940
rect 2430 2905 2470 2910
rect 2430 2885 2445 2905
rect 1165 2865 2445 2885
rect -1000 2840 295 2855
rect -1000 2805 -980 2840
rect -945 2805 295 2840
rect -1000 2790 295 2805
rect 1405 2730 1450 2735
rect 1405 2700 1415 2730
rect 1445 2700 1450 2730
rect 1405 2695 1450 2700
rect 0 2630 295 2685
rect -100 2405 -60 2410
rect -995 2400 -945 2405
rect -100 2400 -95 2405
rect -995 2365 -990 2400
rect -955 2375 -95 2400
rect -65 2375 -60 2405
rect -955 2365 -945 2375
rect -100 2370 -60 2375
rect -995 2360 -945 2365
rect -995 1900 -945 1905
rect -995 1895 -990 1900
rect -1000 1870 -990 1895
rect -995 1865 -990 1870
rect -955 1895 -945 1900
rect -850 1895 -770 1930
rect -115 1900 -75 1905
rect -115 1895 -110 1900
rect -955 1870 -110 1895
rect -80 1870 -75 1900
rect -955 1865 -945 1870
rect -995 1860 -945 1865
rect -850 1850 -770 1870
rect -115 1865 -75 1870
rect 0 1880 50 2630
rect 1405 2590 1425 2695
rect 1360 2585 1450 2590
rect 1360 2575 1415 2585
rect 1360 2490 1385 2575
rect 1410 2555 1415 2575
rect 1445 2555 1450 2585
rect 1410 2550 1450 2555
rect 715 2485 1385 2490
rect 715 2455 720 2485
rect 750 2475 1385 2485
rect 1410 2510 1450 2515
rect 1485 2510 1510 2865
rect 2155 2840 2195 2865
rect 1605 2790 1645 2795
rect 1605 2760 1610 2790
rect 1640 2760 1645 2790
rect 1605 2755 1645 2760
rect 2155 2760 2195 2765
rect 1610 2520 1635 2755
rect 2155 2730 2160 2760
rect 2190 2755 2195 2760
rect 2440 2760 2480 2765
rect 2440 2755 2445 2760
rect 2190 2735 2445 2755
rect 2190 2730 2195 2735
rect 2155 2725 2195 2730
rect 2440 2730 2445 2735
rect 2475 2730 2480 2760
rect 2440 2725 2480 2730
rect 2155 2660 2195 2665
rect 2440 2660 2480 2665
rect 2150 2640 2160 2660
rect 2155 2630 2160 2640
rect 2190 2640 2445 2660
rect 2190 2630 2195 2640
rect 2155 2620 2195 2630
rect 2440 2630 2445 2640
rect 2475 2630 2480 2660
rect 2440 2625 2480 2630
rect 1410 2480 1415 2510
rect 1445 2485 1510 2510
rect 1605 2515 1645 2520
rect 1605 2485 1610 2515
rect 1640 2485 1645 2515
rect 1445 2480 1450 2485
rect 1605 2480 1645 2485
rect 1410 2475 1450 2480
rect 750 2455 755 2475
rect 715 2450 755 2455
rect 200 2410 245 2415
rect 200 2375 205 2410
rect 240 2405 245 2410
rect 880 2405 920 2410
rect 240 2385 885 2405
rect 240 2375 245 2385
rect 200 2370 245 2375
rect 880 2375 885 2385
rect 915 2375 920 2405
rect 880 2370 920 2375
rect 1680 2340 2270 2345
rect 1680 2310 1685 2340
rect 1715 2310 2235 2340
rect 2265 2310 2270 2340
rect 1680 2305 2270 2310
rect 2515 2285 2550 3175
rect 2565 3115 2610 3125
rect 2565 3085 2575 3115
rect 2605 3085 2610 3115
rect 2565 3080 2610 3085
rect 2570 2395 2610 3080
rect 3730 2405 3785 2420
rect 3730 2395 3740 2405
rect 2570 2370 3740 2395
rect 3775 2370 3785 2405
rect 3730 2355 3785 2370
rect 195 2280 665 2285
rect 195 2200 200 2280
rect 230 2200 665 2280
rect 195 2195 665 2200
rect 2015 2225 2550 2285
rect 2015 2195 2390 2225
rect 195 2125 530 2135
rect 195 2045 200 2125
rect 230 2045 530 2125
rect 195 1880 530 2045
rect 0 1790 560 1880
rect 1379 1790 1416 1824
rect 0 0 45 1790
rect 300 1742 320 1790
rect 1361 1766 1407 1772
rect 1361 1742 1366 1766
rect 99 1741 1366 1742
rect 98 1729 1366 1741
rect 1401 1729 1407 1766
rect 98 1723 1407 1729
rect 98 1698 115 1723
rect 86 1658 123 1698
rect 300 1690 320 1723
rect 1361 1721 1407 1723
rect 2350 1630 2390 2195
rect 2575 1950 2615 1960
rect 2575 1920 2580 1950
rect 2610 1945 2615 1950
rect 3555 1945 3640 1970
rect 3730 1955 3785 1970
rect 3730 1945 3740 1955
rect 2610 1925 3740 1945
rect 2610 1920 2615 1925
rect 2575 1910 2615 1920
rect 3555 1885 3640 1925
rect 3730 1920 3740 1925
rect 3775 1920 3785 1955
rect 3730 1905 3785 1920
<< via2 >>
rect -880 5210 -850 5240
rect -105 5210 -75 5240
rect 670 5210 700 5240
rect 1445 5210 1475 5240
rect 2220 5210 2250 5240
rect 2995 5210 3025 5240
rect -980 2805 -945 2840
rect -990 2365 -955 2400
rect -990 1865 -955 1900
rect 3740 2370 3775 2405
rect 3740 1920 3775 1955
<< metal3 >>
rect -885 5240 -825 5245
rect -885 5205 -880 5240
rect -845 5205 -825 5240
rect -110 5240 -50 5245
rect -110 5205 -105 5240
rect -70 5205 -50 5240
rect 665 5240 725 5245
rect 665 5205 670 5240
rect 705 5205 725 5240
rect 1440 5240 1500 5245
rect 1440 5205 1445 5240
rect 1480 5205 1500 5240
rect 2215 5240 2275 5245
rect 2215 5205 2220 5240
rect 2255 5205 2275 5240
rect 2990 5240 3050 5245
rect 2990 5205 2995 5240
rect 3030 5205 3050 5240
rect -900 4310 3710 5165
rect -900 2855 3690 4310
rect -1000 2840 3690 2855
rect -1000 2805 -980 2840
rect -945 2805 3690 2840
rect -1000 2790 3690 2805
rect -1000 2400 -945 2415
rect -1000 2365 -990 2400
rect -955 2365 -945 2400
rect -1000 2350 -945 2365
rect -1000 1900 -945 1915
rect -1000 1865 -990 1900
rect -955 1865 -945 1900
rect -1000 1850 -945 1865
rect -900 -180 3690 2790
rect 3730 2405 3785 2420
rect 3730 2370 3740 2405
rect 3775 2370 3785 2405
rect 3730 2355 3785 2370
rect 3730 1955 3785 1970
rect 3730 1920 3740 1955
rect 3775 1920 3785 1955
rect 3730 1905 3785 1920
rect -890 -210 3690 -180
<< via3 >>
rect -880 5210 -850 5240
rect -850 5210 -845 5240
rect -880 5205 -845 5210
rect -105 5210 -75 5240
rect -75 5210 -70 5240
rect -105 5205 -70 5210
rect 670 5210 700 5240
rect 700 5210 705 5240
rect 670 5205 705 5210
rect 1445 5210 1475 5240
rect 1475 5210 1480 5240
rect 1445 5205 1480 5210
rect 2220 5210 2250 5240
rect 2250 5210 2255 5240
rect 2220 5205 2255 5210
rect 2995 5210 3025 5240
rect 3025 5210 3030 5240
rect 2995 5205 3030 5210
rect -990 2365 -955 2400
rect -990 1865 -955 1900
rect 3740 2370 3775 2405
rect 3740 1920 3775 1955
<< mimcap >>
rect -885 5120 -195 5145
rect -885 5035 -860 5120
rect -775 5035 -195 5120
rect -885 4455 -195 5035
rect -110 5120 580 5145
rect -110 5035 -85 5120
rect 0 5035 580 5120
rect -110 4455 580 5035
rect 665 5120 1355 5145
rect 665 5035 690 5120
rect 775 5035 1355 5120
rect 665 4455 1355 5035
rect 1440 5120 2130 5145
rect 1440 5035 1465 5120
rect 1550 5035 2130 5120
rect 1440 4455 2130 5035
rect 2215 5120 2905 5145
rect 2215 5035 2240 5120
rect 2325 5035 2905 5120
rect 2215 4455 2905 5035
rect 2990 5120 3680 5145
rect 2990 5035 3015 5120
rect 3100 5035 3680 5120
rect 2990 4455 3680 5035
rect -870 2430 1350 4370
rect -870 2350 -850 2430
rect -770 2350 1350 2430
rect -870 2150 1350 2350
rect 1440 2420 3660 4370
rect 1440 2340 3550 2420
rect 3630 2340 3660 2420
rect 1440 2150 3660 2340
rect -870 1930 1350 2060
rect -870 1850 -850 1930
rect -770 1850 1350 1930
rect -870 -160 1350 1850
rect 1440 1970 3660 2060
rect 1440 1890 3550 1970
rect 3630 1890 3660 1970
rect 1440 -160 3660 1890
<< mimcapcontact >>
rect -860 5035 -775 5120
rect -85 5035 0 5120
rect 690 5035 775 5120
rect 1465 5035 1550 5120
rect 2240 5035 2325 5120
rect 3015 5035 3100 5120
rect -850 2350 -770 2430
rect 3550 2340 3630 2420
rect -850 1850 -770 1930
rect 3550 1890 3630 1970
<< metal4 >>
rect -885 5240 -825 5245
rect -885 5205 -880 5240
rect -845 5205 -825 5240
rect -885 5145 -825 5205
rect -110 5240 -50 5245
rect -110 5205 -105 5240
rect -70 5205 -50 5240
rect -110 5145 -50 5205
rect 665 5240 725 5245
rect 665 5205 670 5240
rect 705 5205 725 5240
rect 665 5145 725 5205
rect 1440 5240 1500 5245
rect 1440 5205 1445 5240
rect 1480 5205 1500 5240
rect 1440 5145 1500 5205
rect 2215 5240 2275 5245
rect 2215 5205 2220 5240
rect 2255 5205 2275 5240
rect 2215 5145 2275 5205
rect 2990 5240 3050 5245
rect 2990 5205 2995 5240
rect 3030 5205 3050 5240
rect 2990 5145 3050 5205
rect -885 5120 -755 5145
rect -885 5035 -860 5120
rect -775 5035 -755 5120
rect -885 5025 -755 5035
rect -110 5120 20 5145
rect -110 5035 -85 5120
rect 0 5035 20 5120
rect -110 5025 20 5035
rect 665 5120 795 5145
rect 665 5035 690 5120
rect 775 5035 795 5120
rect 665 5025 795 5035
rect 1440 5120 1570 5145
rect 1440 5035 1465 5120
rect 1550 5035 1570 5120
rect 1440 5025 1570 5035
rect 2215 5120 2345 5145
rect 2215 5035 2240 5120
rect 2325 5035 2345 5120
rect 2215 5025 2345 5035
rect 2990 5120 3120 5145
rect 2990 5035 3015 5120
rect 3100 5035 3120 5120
rect 2990 5025 3120 5035
rect -1000 2430 -745 2440
rect -1000 2400 -850 2430
rect -1000 2365 -990 2400
rect -955 2365 -850 2400
rect -1000 2350 -850 2365
rect -770 2350 -745 2430
rect -1000 2325 -745 2350
rect 3520 2420 3790 2440
rect 3520 2340 3550 2420
rect 3630 2405 3790 2420
rect 3630 2370 3740 2405
rect 3775 2370 3790 2405
rect 3630 2340 3790 2370
rect 3520 2320 3790 2340
rect 3525 1970 3795 1990
rect -1000 1930 -745 1945
rect -1000 1900 -850 1930
rect -1000 1865 -990 1900
rect -955 1865 -850 1900
rect -1000 1850 -850 1865
rect -770 1850 -745 1930
rect 3525 1890 3550 1970
rect 3630 1955 3795 1970
rect 3630 1920 3740 1955
rect 3775 1920 3795 1955
rect 3630 1890 3795 1920
rect 3525 1870 3795 1890
rect -1000 1830 -745 1850
use bias_cg  bias_cg_0 ~/Documents/Final/bi-directional-A-D-A-converter/layout
timestamp 1702648396
transform 1 0 385 0 1 970
box -385 -970 2311 660
use com_di  com_di_0 ~/Documents/Final/bi-directional-A-D-A-converter/layout
timestamp 1702662166
transform 1 0 1085 0 1 2870
box -855 -395 1330 635
use middle  middle_0 ~/Documents/Final/bi-directional-A-D-A-converter/layout
timestamp 1702643716
transform 1 0 270 0 1 2060
box 50 -410 2085 405
<< labels >>
rlabel metal1 -1000 2755 -1000 2755 1 RST
port 4 n
rlabel metal1 3725 2745 3725 2745 1 SEN
port 5 n
rlabel metal1 -1000 1985 -1000 1985 1 PRE
port 6 n
rlabel metal1 -1000 2545 -1000 2545 1 ENAD
port 7 n
rlabel metal1 -1000 1678 -1000 1678 1 SH
port 8 n
rlabel metal1 -1003 2145 -1003 2145 1 Vref-
port 9 n
rlabel metal1 3746 2234 3746 2234 1 Vref+
port 10 n
rlabel metal1 3725 2645 3725 2645 1 D
port 11 n
<< end >>
