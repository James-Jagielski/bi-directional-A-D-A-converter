magic
tech sky130A
timestamp 1702614174
<< nwell >>
rect 1051 125 1400 126
rect -270 -20 2199 125
rect 825 -21 1400 -20
rect 825 -175 1063 -21
<< nmos >>
rect -60 -190 -45 -90
rect 85 -190 100 -90
rect 150 -190 165 -90
rect 295 -190 310 -90
rect 440 -190 455 -90
rect 505 -190 520 -90
rect 650 -190 665 -90
rect 1340 -190 1355 -90
rect 1485 -190 1500 -90
rect 1550 -190 1565 -90
rect 1695 -190 1710 -90
rect 1840 -190 1855 -90
rect 1905 -190 1920 -90
rect 2050 -190 2065 -90
rect -125 -385 -110 -285
rect -60 -385 -45 -285
rect 5 -385 20 -285
rect 195 -385 210 -285
rect 260 -385 275 -285
rect 330 -385 345 -285
rect 395 -385 410 -285
rect 585 -385 600 -285
rect 650 -385 665 -285
rect 715 -385 730 -285
rect 940 -310 955 -210
rect 940 -440 955 -340
rect 1275 -385 1290 -285
rect 1340 -385 1355 -285
rect 1405 -385 1420 -285
rect 1595 -385 1610 -285
rect 1660 -385 1675 -285
rect 1730 -385 1745 -285
rect 1795 -385 1810 -285
rect 1985 -385 2000 -285
rect 2050 -385 2065 -285
rect 2115 -385 2130 -285
<< pmos >>
rect -105 0 -90 100
rect -40 0 -25 100
rect 25 0 40 100
rect 90 0 105 100
rect 155 0 170 100
rect 220 0 235 100
rect 370 0 385 100
rect 435 0 450 100
rect 500 0 515 100
rect 565 0 580 100
rect 630 0 645 100
rect 695 0 710 100
rect 940 0 955 100
rect 1295 0 1310 100
rect 1360 0 1375 100
rect 1425 0 1440 100
rect 1490 0 1505 100
rect 1555 0 1570 100
rect 1620 0 1635 100
rect 940 -155 955 -55
rect 1770 0 1785 100
rect 1835 0 1850 100
rect 1900 0 1915 100
rect 1965 0 1980 100
rect 2030 0 2045 100
rect 2095 0 2110 100
<< ndiff >>
rect -110 -105 -60 -90
rect -110 -175 -95 -105
rect -75 -175 -60 -105
rect -110 -190 -60 -175
rect -45 -105 5 -90
rect -45 -175 -30 -105
rect -10 -175 5 -105
rect -45 -190 5 -175
rect 35 -105 85 -90
rect 35 -175 50 -105
rect 70 -175 85 -105
rect 35 -190 85 -175
rect 100 -105 150 -90
rect 100 -175 115 -105
rect 135 -175 150 -105
rect 100 -190 150 -175
rect 165 -105 215 -90
rect 165 -175 180 -105
rect 200 -175 215 -105
rect 165 -190 215 -175
rect 245 -105 295 -90
rect 245 -175 260 -105
rect 280 -175 295 -105
rect 245 -190 295 -175
rect 310 -105 360 -90
rect 310 -175 325 -105
rect 345 -175 360 -105
rect 310 -190 360 -175
rect 390 -105 440 -90
rect 390 -175 405 -105
rect 425 -175 440 -105
rect 390 -190 440 -175
rect 455 -105 505 -90
rect 455 -175 470 -105
rect 490 -175 505 -105
rect 455 -190 505 -175
rect 520 -105 570 -90
rect 520 -175 535 -105
rect 555 -175 570 -105
rect 520 -190 570 -175
rect 600 -105 650 -90
rect 600 -175 615 -105
rect 635 -175 650 -105
rect 600 -190 650 -175
rect 665 -105 715 -90
rect 665 -175 680 -105
rect 700 -175 715 -105
rect 1290 -105 1340 -90
rect 665 -190 715 -175
rect 1290 -175 1305 -105
rect 1325 -175 1340 -105
rect 1290 -190 1340 -175
rect 1355 -105 1405 -90
rect 1355 -175 1370 -105
rect 1390 -175 1405 -105
rect 1355 -190 1405 -175
rect 1435 -105 1485 -90
rect 1435 -175 1450 -105
rect 1470 -175 1485 -105
rect 1435 -190 1485 -175
rect 1500 -105 1550 -90
rect 1500 -175 1515 -105
rect 1535 -175 1550 -105
rect 1500 -190 1550 -175
rect 1565 -105 1615 -90
rect 1565 -175 1580 -105
rect 1600 -175 1615 -105
rect 1565 -190 1615 -175
rect 1645 -105 1695 -90
rect 1645 -175 1660 -105
rect 1680 -175 1695 -105
rect 1645 -190 1695 -175
rect 1710 -105 1760 -90
rect 1710 -175 1725 -105
rect 1745 -175 1760 -105
rect 1710 -190 1760 -175
rect 1790 -105 1840 -90
rect 1790 -175 1805 -105
rect 1825 -175 1840 -105
rect 1790 -190 1840 -175
rect 1855 -105 1905 -90
rect 1855 -175 1870 -105
rect 1890 -175 1905 -105
rect 1855 -190 1905 -175
rect 1920 -105 1970 -90
rect 1920 -175 1935 -105
rect 1955 -175 1970 -105
rect 1920 -190 1970 -175
rect 2000 -105 2050 -90
rect 2000 -175 2015 -105
rect 2035 -175 2050 -105
rect 2000 -190 2050 -175
rect 2065 -105 2115 -90
rect 2065 -175 2080 -105
rect 2100 -175 2115 -105
rect 2065 -190 2115 -175
rect 890 -225 940 -210
rect -175 -300 -125 -285
rect -175 -370 -160 -300
rect -140 -370 -125 -300
rect -175 -385 -125 -370
rect -110 -300 -60 -285
rect -110 -370 -95 -300
rect -75 -370 -60 -300
rect -110 -385 -60 -370
rect -45 -300 5 -285
rect -45 -370 -30 -300
rect -10 -370 5 -300
rect -45 -385 5 -370
rect 20 -300 70 -285
rect 20 -370 35 -300
rect 55 -370 70 -300
rect 20 -385 70 -370
rect 145 -300 195 -285
rect 145 -370 160 -300
rect 180 -370 195 -300
rect 145 -385 195 -370
rect 210 -300 260 -285
rect 210 -370 225 -300
rect 245 -370 260 -300
rect 210 -385 260 -370
rect 275 -300 330 -285
rect 275 -370 290 -300
rect 315 -370 330 -300
rect 275 -385 330 -370
rect 345 -300 395 -285
rect 345 -370 360 -300
rect 380 -370 395 -300
rect 345 -385 395 -370
rect 410 -300 460 -285
rect 410 -370 425 -300
rect 445 -370 460 -300
rect 410 -385 460 -370
rect 535 -300 585 -285
rect 535 -370 550 -300
rect 570 -370 585 -300
rect 535 -385 585 -370
rect 600 -300 650 -285
rect 600 -370 615 -300
rect 635 -370 650 -300
rect 600 -385 650 -370
rect 665 -300 715 -285
rect 665 -370 680 -300
rect 700 -370 715 -300
rect 665 -385 715 -370
rect 730 -300 780 -285
rect 730 -370 745 -300
rect 765 -370 780 -300
rect 890 -295 905 -225
rect 925 -295 940 -225
rect 890 -310 940 -295
rect 955 -225 1005 -210
rect 955 -295 969 -225
rect 990 -295 1005 -225
rect 955 -310 1005 -295
rect 730 -385 780 -370
rect 890 -356 940 -340
rect 890 -427 905 -356
rect 926 -427 940 -356
rect 890 -440 940 -427
rect 955 -356 1005 -340
rect 955 -427 967 -356
rect 988 -427 1005 -356
rect 1225 -300 1275 -285
rect 1225 -370 1240 -300
rect 1260 -370 1275 -300
rect 1225 -385 1275 -370
rect 1290 -300 1340 -285
rect 1290 -370 1305 -300
rect 1325 -370 1340 -300
rect 1290 -385 1340 -370
rect 1355 -300 1405 -285
rect 1355 -370 1370 -300
rect 1390 -370 1405 -300
rect 1355 -385 1405 -370
rect 1420 -300 1470 -285
rect 1420 -370 1435 -300
rect 1455 -370 1470 -300
rect 1420 -385 1470 -370
rect 1545 -300 1595 -285
rect 1545 -370 1560 -300
rect 1580 -370 1595 -300
rect 1545 -385 1595 -370
rect 1610 -300 1660 -285
rect 1610 -370 1625 -300
rect 1645 -370 1660 -300
rect 1610 -385 1660 -370
rect 1675 -300 1730 -285
rect 1675 -370 1690 -300
rect 1715 -370 1730 -300
rect 1675 -385 1730 -370
rect 1745 -300 1795 -285
rect 1745 -370 1760 -300
rect 1780 -370 1795 -300
rect 1745 -385 1795 -370
rect 1810 -300 1860 -285
rect 1810 -370 1825 -300
rect 1845 -370 1860 -300
rect 1810 -385 1860 -370
rect 1935 -300 1985 -285
rect 1935 -370 1950 -300
rect 1970 -370 1985 -300
rect 1935 -385 1985 -370
rect 2000 -300 2050 -285
rect 2000 -370 2015 -300
rect 2035 -370 2050 -300
rect 2000 -385 2050 -370
rect 2065 -300 2115 -285
rect 2065 -370 2080 -300
rect 2100 -370 2115 -300
rect 2065 -385 2115 -370
rect 2130 -300 2180 -285
rect 2130 -370 2145 -300
rect 2165 -370 2180 -300
rect 2130 -385 2180 -370
rect 955 -440 1005 -427
<< pdiff >>
rect -155 85 -105 100
rect -155 15 -140 85
rect -120 15 -105 85
rect -155 0 -105 15
rect -90 85 -40 100
rect -90 15 -75 85
rect -55 15 -40 85
rect -90 0 -40 15
rect -25 85 25 100
rect -25 15 -10 85
rect 10 15 25 85
rect -25 0 25 15
rect 40 85 90 100
rect 40 15 55 85
rect 75 15 90 85
rect 40 0 90 15
rect 105 0 155 100
rect 170 85 220 100
rect 170 15 185 85
rect 205 15 220 85
rect 170 0 220 15
rect 235 85 285 100
rect 235 15 250 85
rect 270 15 285 85
rect 235 0 285 15
rect 320 85 370 100
rect 320 15 335 85
rect 355 15 370 85
rect 320 0 370 15
rect 385 85 435 100
rect 385 15 400 85
rect 420 15 435 85
rect 385 0 435 15
rect 450 0 500 100
rect 515 85 565 100
rect 515 15 530 85
rect 550 15 565 85
rect 515 0 565 15
rect 580 85 630 100
rect 580 15 595 85
rect 615 15 630 85
rect 580 0 630 15
rect 645 85 695 100
rect 645 15 660 85
rect 680 15 695 85
rect 645 0 695 15
rect 710 85 760 100
rect 710 15 725 85
rect 745 15 760 85
rect 890 84 940 100
rect 710 0 760 15
rect 890 13 906 84
rect 927 13 940 84
rect 890 0 940 13
rect 955 86 1005 100
rect 955 15 968 86
rect 989 15 1005 86
rect 955 0 1005 15
rect 1245 85 1295 100
rect 1245 15 1260 85
rect 1280 15 1295 85
rect 1245 0 1295 15
rect 1310 85 1360 100
rect 1310 15 1325 85
rect 1345 15 1360 85
rect 1310 0 1360 15
rect 1375 85 1425 100
rect 1375 15 1390 85
rect 1410 15 1425 85
rect 1375 0 1425 15
rect 1440 85 1490 100
rect 1440 15 1455 85
rect 1475 15 1490 85
rect 1440 0 1490 15
rect 1505 0 1555 100
rect 1570 85 1620 100
rect 1570 15 1585 85
rect 1605 15 1620 85
rect 1570 0 1620 15
rect 1635 85 1685 100
rect 1635 15 1650 85
rect 1670 15 1685 85
rect 1635 0 1685 15
rect 890 -70 940 -55
rect 890 -140 905 -70
rect 925 -140 940 -70
rect 890 -155 940 -140
rect 955 -70 1005 -55
rect 955 -140 970 -70
rect 990 -140 1005 -70
rect 1720 85 1770 100
rect 1720 15 1735 85
rect 1755 15 1770 85
rect 1720 0 1770 15
rect 1785 85 1835 100
rect 1785 15 1800 85
rect 1820 15 1835 85
rect 1785 0 1835 15
rect 1850 0 1900 100
rect 1915 85 1965 100
rect 1915 15 1930 85
rect 1950 15 1965 85
rect 1915 0 1965 15
rect 1980 85 2030 100
rect 1980 15 1995 85
rect 2015 15 2030 85
rect 1980 0 2030 15
rect 2045 85 2095 100
rect 2045 15 2060 85
rect 2080 15 2095 85
rect 2045 0 2095 15
rect 2110 85 2160 100
rect 2110 15 2125 85
rect 2145 15 2160 85
rect 2110 0 2160 15
rect 955 -155 1005 -140
<< ndiffc >>
rect -95 -175 -75 -105
rect -30 -175 -10 -105
rect 50 -175 70 -105
rect 115 -175 135 -105
rect 180 -175 200 -105
rect 260 -175 280 -105
rect 325 -175 345 -105
rect 405 -175 425 -105
rect 470 -175 490 -105
rect 535 -175 555 -105
rect 615 -175 635 -105
rect 680 -175 700 -105
rect 1305 -175 1325 -105
rect 1370 -175 1390 -105
rect 1450 -175 1470 -105
rect 1515 -175 1535 -105
rect 1580 -175 1600 -105
rect 1660 -175 1680 -105
rect 1725 -175 1745 -105
rect 1805 -175 1825 -105
rect 1870 -175 1890 -105
rect 1935 -175 1955 -105
rect 2015 -175 2035 -105
rect 2080 -175 2100 -105
rect -160 -370 -140 -300
rect -95 -370 -75 -300
rect -30 -370 -10 -300
rect 35 -370 55 -300
rect 160 -370 180 -300
rect 225 -370 245 -300
rect 290 -370 315 -300
rect 360 -370 380 -300
rect 425 -370 445 -300
rect 550 -370 570 -300
rect 615 -370 635 -300
rect 680 -370 700 -300
rect 745 -370 765 -300
rect 905 -295 925 -225
rect 969 -295 990 -225
rect 905 -427 926 -356
rect 967 -427 988 -356
rect 1240 -370 1260 -300
rect 1305 -370 1325 -300
rect 1370 -370 1390 -300
rect 1435 -370 1455 -300
rect 1560 -370 1580 -300
rect 1625 -370 1645 -300
rect 1690 -370 1715 -300
rect 1760 -370 1780 -300
rect 1825 -370 1845 -300
rect 1950 -370 1970 -300
rect 2015 -370 2035 -300
rect 2080 -370 2100 -300
rect 2145 -370 2165 -300
<< pdiffc >>
rect -140 15 -120 85
rect -75 15 -55 85
rect -10 15 10 85
rect 55 15 75 85
rect 185 15 205 85
rect 250 15 270 85
rect 335 15 355 85
rect 400 15 420 85
rect 530 15 550 85
rect 595 15 615 85
rect 660 15 680 85
rect 725 15 745 85
rect 906 13 927 84
rect 968 15 989 86
rect 1260 15 1280 85
rect 1325 15 1345 85
rect 1390 15 1410 85
rect 1455 15 1475 85
rect 1585 15 1605 85
rect 1650 15 1670 85
rect 905 -140 925 -70
rect 970 -140 990 -70
rect 1735 15 1755 85
rect 1800 15 1820 85
rect 1930 15 1950 85
rect 1995 15 2015 85
rect 2060 15 2080 85
rect 2125 15 2145 85
<< psubdiff >>
rect -255 -300 -205 -285
rect -255 -370 -240 -300
rect -220 -370 -205 -300
rect -255 -385 -205 -370
rect 1145 -300 1195 -285
rect 1145 -370 1160 -300
rect 1180 -370 1195 -300
rect 1145 -385 1195 -370
<< nsubdiff >>
rect -250 85 -200 100
rect -250 15 -235 85
rect -215 15 -200 85
rect -250 0 -200 15
rect 1150 85 1200 100
rect 1150 15 1165 85
rect 1185 15 1200 85
rect 1150 0 1200 15
<< psubdiffcont >>
rect -240 -370 -220 -300
rect 1160 -370 1180 -300
<< nsubdiffcont >>
rect -235 15 -215 85
rect 1165 15 1185 85
<< poly >>
rect -188 205 -146 214
rect -188 180 -179 205
rect -156 180 -146 205
rect -188 170 -146 180
rect -117 204 -76 213
rect -117 180 -108 204
rect -84 180 -76 204
rect 694 206 733 214
rect -117 171 -76 180
rect 25 183 647 199
rect 694 183 702 206
rect 724 183 733 206
rect 25 182 645 183
rect -188 -36 -172 170
rect -105 100 -90 171
rect -40 100 -25 165
rect 25 115 41 182
rect 175 150 215 160
rect 175 130 185 150
rect 205 130 215 150
rect 390 150 430 160
rect 175 125 215 130
rect 25 100 40 115
rect 90 100 105 125
rect 155 110 235 125
rect 155 100 170 110
rect 220 100 235 110
rect -105 -15 -90 0
rect -40 -36 -25 0
rect 25 -15 40 0
rect 90 -15 105 0
rect 155 -15 170 0
rect 220 -15 235 0
rect -188 -51 -25 -36
rect 85 -47 120 -40
rect 85 -66 93 -47
rect 112 -66 120 -47
rect 85 -75 120 -66
rect -60 -90 -45 -75
rect 85 -90 100 -75
rect 150 -90 165 -75
rect 295 -90 310 145
rect 390 130 400 150
rect 420 130 430 150
rect 390 125 430 130
rect 553 144 592 156
rect 370 110 450 125
rect 553 124 563 144
rect 583 124 592 144
rect 370 100 385 110
rect 435 100 450 110
rect 500 100 515 115
rect 553 114 592 124
rect 565 100 580 114
rect 630 100 645 182
rect 694 173 733 183
rect 1212 205 1254 214
rect 1212 180 1221 205
rect 1244 180 1254 205
rect 694 113 710 173
rect 1212 170 1254 180
rect 1283 204 1324 213
rect 1283 180 1292 204
rect 1316 180 1324 204
rect 2094 206 2133 214
rect 1283 171 1324 180
rect 1425 183 2047 199
rect 2094 183 2102 206
rect 2124 183 2133 206
rect 1425 182 2045 183
rect 856 116 955 125
rect 695 100 710 113
rect 840 110 955 116
rect 840 108 872 110
rect 840 91 848 108
rect 865 91 872 108
rect 940 100 955 110
rect 840 83 872 91
rect 370 -15 385 0
rect 435 -15 450 0
rect 500 -15 515 0
rect 565 -15 580 0
rect 630 -15 645 0
rect 695 -15 710 0
rect 940 -15 955 0
rect 1212 -36 1228 170
rect 1295 100 1310 171
rect 1360 100 1375 165
rect 1425 115 1441 182
rect 1575 150 1615 160
rect 1575 130 1585 150
rect 1605 130 1615 150
rect 1790 150 1830 160
rect 1575 125 1615 130
rect 1425 100 1440 115
rect 1490 100 1505 125
rect 1555 110 1635 125
rect 1555 100 1570 110
rect 1620 100 1635 110
rect 1295 -15 1310 0
rect 1360 -36 1375 0
rect 1425 -15 1440 0
rect 1490 -15 1505 0
rect 1555 -15 1570 0
rect 1620 -15 1635 0
rect 485 -48 520 -40
rect 485 -67 493 -48
rect 512 -67 520 -48
rect 940 -55 955 -40
rect 1212 -51 1375 -36
rect 1485 -47 1520 -40
rect 485 -75 520 -67
rect 440 -90 455 -75
rect 505 -90 520 -75
rect 650 -90 665 -75
rect 1485 -66 1493 -47
rect 1512 -66 1520 -47
rect 1485 -75 1520 -66
rect 1340 -90 1355 -75
rect 1485 -90 1500 -75
rect 1550 -90 1565 -75
rect 1695 -90 1710 145
rect 1790 130 1800 150
rect 1820 130 1830 150
rect 1790 125 1830 130
rect 1953 144 1992 156
rect 1770 110 1850 125
rect 1953 124 1963 144
rect 1983 124 1992 144
rect 1770 100 1785 110
rect 1835 100 1850 110
rect 1900 100 1915 115
rect 1953 114 1992 124
rect 1965 100 1980 114
rect 2030 100 2045 182
rect 2094 173 2133 183
rect 2094 113 2110 173
rect 2095 100 2110 113
rect 1770 -15 1785 0
rect 1835 -15 1850 0
rect 1900 -15 1915 0
rect 1965 -15 1980 0
rect 2030 -15 2045 0
rect 2095 -15 2110 0
rect 1885 -48 1920 -40
rect 1885 -67 1893 -48
rect 1912 -67 1920 -48
rect 1885 -75 1920 -67
rect 1840 -90 1855 -75
rect 1905 -90 1920 -75
rect 2050 -90 2065 -75
rect -60 -205 -45 -190
rect 85 -205 100 -190
rect 150 -200 165 -190
rect -85 -215 -45 -205
rect 150 -215 210 -200
rect 295 -205 310 -190
rect 440 -200 455 -190
rect -85 -235 -75 -215
rect -55 -235 -45 -215
rect -85 -245 -45 -235
rect -125 -285 -110 -270
rect -60 -285 -45 -270
rect 5 -285 20 -270
rect 195 -285 210 -215
rect 395 -215 455 -200
rect 505 -205 520 -190
rect 650 -205 665 -190
rect 650 -215 690 -205
rect 940 -210 955 -155
rect 1340 -205 1355 -190
rect 1485 -205 1500 -190
rect 1550 -200 1565 -190
rect 260 -285 275 -270
rect 330 -285 345 -270
rect 395 -285 410 -215
rect 650 -235 660 -215
rect 680 -235 690 -215
rect 650 -245 690 -235
rect 585 -285 600 -270
rect 650 -285 665 -270
rect 715 -285 730 -270
rect 1315 -215 1355 -205
rect 1550 -215 1610 -200
rect 1695 -205 1710 -190
rect 1840 -200 1855 -190
rect 1315 -235 1325 -215
rect 1345 -235 1355 -215
rect 1315 -245 1355 -235
rect 1275 -285 1290 -270
rect 1340 -285 1355 -270
rect 1405 -285 1420 -270
rect 1595 -285 1610 -215
rect 1795 -215 1855 -200
rect 1905 -205 1920 -190
rect 2050 -205 2065 -190
rect 2050 -215 2090 -205
rect 1660 -285 1675 -270
rect 1730 -285 1745 -270
rect 1795 -285 1810 -215
rect 2050 -235 2060 -215
rect 2080 -235 2090 -215
rect 2050 -245 2090 -235
rect 1985 -285 2000 -270
rect 2050 -285 2065 -270
rect 2115 -285 2130 -270
rect 940 -340 955 -310
rect -125 -455 -110 -385
rect -60 -398 -45 -385
rect -77 -407 -41 -398
rect -77 -427 -69 -407
rect -50 -427 -41 -407
rect 5 -420 20 -385
rect -77 -434 -41 -427
rect -137 -463 -99 -455
rect -137 -485 -128 -463
rect -107 -485 -99 -463
rect 4 -464 21 -420
rect 195 -425 210 -385
rect 260 -400 275 -385
rect 330 -400 345 -385
rect 395 -425 410 -385
rect 585 -399 600 -385
rect 195 -440 410 -425
rect 568 -407 604 -399
rect 568 -427 577 -407
rect 596 -427 604 -407
rect 568 -435 604 -427
rect 650 -464 665 -385
rect 715 -455 730 -385
rect 4 -480 665 -464
rect 701 -464 740 -455
rect -137 -494 -99 -485
rect 701 -486 710 -464
rect 731 -486 740 -464
rect 940 -465 955 -440
rect 1275 -455 1290 -385
rect 1340 -398 1355 -385
rect 1323 -407 1359 -398
rect 1323 -427 1331 -407
rect 1350 -427 1359 -407
rect 1405 -420 1420 -385
rect 1323 -434 1359 -427
rect 1263 -463 1301 -455
rect 701 -494 740 -486
rect 1263 -485 1272 -463
rect 1293 -485 1301 -463
rect 1404 -464 1421 -420
rect 1595 -425 1610 -385
rect 1660 -400 1675 -385
rect 1730 -400 1745 -385
rect 1795 -425 1810 -385
rect 1985 -399 2000 -385
rect 1595 -440 1810 -425
rect 1968 -407 2004 -399
rect 1968 -427 1977 -407
rect 1996 -427 2004 -407
rect 1968 -435 2004 -427
rect 2050 -464 2065 -385
rect 2115 -455 2130 -385
rect 1404 -480 2065 -464
rect 2101 -464 2140 -455
rect 1263 -494 1301 -485
rect 2101 -486 2110 -464
rect 2131 -486 2140 -464
rect 2101 -494 2140 -486
<< polycont >>
rect -179 180 -156 205
rect -108 180 -84 204
rect 702 183 724 206
rect 185 130 205 150
rect 93 -66 112 -47
rect 400 130 420 150
rect 563 124 583 144
rect 1221 180 1244 205
rect 1292 180 1316 204
rect 2102 183 2124 206
rect 848 91 865 108
rect 1585 130 1605 150
rect 493 -67 512 -48
rect 1493 -66 1512 -47
rect 1800 130 1820 150
rect 1963 124 1983 144
rect 1893 -67 1912 -48
rect -75 -235 -55 -215
rect 660 -235 680 -215
rect 1325 -235 1345 -215
rect 2060 -235 2080 -215
rect -69 -427 -50 -407
rect -128 -485 -107 -463
rect 577 -427 596 -407
rect 710 -486 731 -464
rect 1331 -427 1350 -407
rect 1272 -485 1293 -463
rect 1977 -427 1996 -407
rect 2110 -486 2131 -464
<< locali >>
rect -188 205 -146 214
rect -188 180 -179 205
rect -156 180 -146 205
rect -188 170 -146 180
rect -117 204 -76 213
rect 694 206 733 215
rect 694 204 702 206
rect -117 180 -108 204
rect -84 183 702 204
rect 724 183 733 206
rect -84 180 733 183
rect -117 179 733 180
rect -117 171 -76 179
rect 694 173 733 179
rect 1212 205 1254 214
rect 1212 180 1221 205
rect 1244 180 1254 205
rect 1212 170 1254 180
rect 1283 204 1324 213
rect 2094 206 2133 215
rect 2094 204 2102 206
rect 1283 180 1292 204
rect 1316 183 2102 204
rect 2124 183 2133 206
rect 1316 180 2133 183
rect 1283 179 2133 180
rect 1283 171 1324 179
rect 2094 173 2133 179
rect 175 150 215 160
rect 175 130 185 150
rect 205 130 215 150
rect 175 120 215 130
rect 390 150 430 160
rect 390 130 400 150
rect 420 130 430 150
rect 390 120 430 130
rect 553 144 592 156
rect 553 124 563 144
rect 583 124 592 144
rect 553 114 592 124
rect 670 134 920 154
rect 670 95 689 134
rect 840 108 872 116
rect -245 85 -205 95
rect -245 15 -235 85
rect -215 15 -205 85
rect -150 85 -110 95
rect -150 25 -140 85
rect -245 5 -205 15
rect -185 15 -140 25
rect -120 15 -110 85
rect -185 5 -110 15
rect -85 85 20 95
rect -85 15 -75 85
rect -55 15 -10 85
rect 10 15 20 85
rect -85 5 20 15
rect 45 85 85 95
rect 45 15 55 85
rect 75 15 85 85
rect 45 5 85 15
rect 175 85 215 95
rect 175 15 185 85
rect 205 15 215 85
rect 175 5 215 15
rect 240 85 280 95
rect 240 15 250 85
rect 270 15 280 85
rect 240 5 280 15
rect 325 85 365 95
rect 325 15 335 85
rect 355 15 365 85
rect 325 5 365 15
rect 390 85 430 95
rect 390 15 400 85
rect 420 15 430 85
rect 390 5 430 15
rect 520 85 560 95
rect 520 15 530 85
rect 550 15 560 85
rect 520 5 560 15
rect 585 85 690 95
rect 585 15 595 85
rect 615 15 660 85
rect 680 15 690 85
rect 585 5 690 15
rect 715 85 755 95
rect 715 15 725 85
rect 745 25 755 85
rect 840 91 848 108
rect 865 91 872 108
rect 900 96 920 134
rect 1025 133 1337 153
rect 1025 97 1046 133
rect 840 83 872 91
rect 894 84 937 96
rect 745 15 790 25
rect 715 5 790 15
rect -185 -255 -165 5
rect -85 -15 -65 5
rect -145 -35 -65 -15
rect 670 -15 690 5
rect 670 -35 750 -15
rect -145 -205 -125 -35
rect 85 -47 520 -40
rect 85 -66 93 -47
rect 112 -48 520 -47
rect 112 -60 493 -48
rect 112 -66 120 -60
rect 85 -75 120 -66
rect 190 -95 210 -60
rect 395 -95 415 -60
rect 485 -67 493 -60
rect 512 -67 520 -48
rect 485 -75 520 -67
rect -105 -105 -65 -95
rect -105 -175 -95 -105
rect -75 -175 -65 -105
rect -105 -185 -65 -175
rect -40 -105 0 -95
rect -40 -175 -30 -105
rect -10 -175 0 -105
rect -40 -185 0 -175
rect 40 -105 80 -95
rect 40 -175 50 -105
rect 70 -175 80 -105
rect 40 -185 80 -175
rect 105 -105 145 -95
rect 105 -175 115 -105
rect 135 -175 145 -105
rect 105 -185 145 -175
rect 170 -105 210 -95
rect 170 -175 180 -105
rect 200 -175 210 -105
rect 170 -185 210 -175
rect 250 -105 290 -95
rect 250 -175 260 -105
rect 280 -175 290 -105
rect 250 -185 290 -175
rect 315 -105 355 -95
rect 315 -175 325 -105
rect 345 -175 355 -105
rect 315 -185 355 -175
rect 395 -105 435 -95
rect 395 -175 405 -105
rect 425 -175 435 -105
rect 395 -185 435 -175
rect 460 -105 500 -95
rect 460 -175 470 -105
rect 490 -175 500 -105
rect 460 -185 500 -175
rect 525 -105 565 -95
rect 525 -175 535 -105
rect 555 -175 565 -105
rect 525 -185 565 -175
rect 605 -105 645 -95
rect 605 -175 615 -105
rect 635 -175 645 -105
rect 605 -185 645 -175
rect 670 -105 710 -95
rect 670 -175 680 -105
rect 700 -175 710 -105
rect 670 -185 710 -175
rect -20 -205 0 -185
rect 335 -205 355 -185
rect 605 -205 625 -185
rect 730 -205 750 -35
rect -145 -215 -45 -205
rect -145 -225 -75 -215
rect -85 -235 -75 -225
rect -55 -235 -45 -215
rect -20 -225 625 -205
rect 650 -215 750 -205
rect -85 -245 -45 -235
rect 650 -235 660 -215
rect 680 -225 750 -215
rect 680 -235 690 -225
rect 650 -245 690 -235
rect -185 -275 -150 -255
rect -170 -290 -150 -275
rect -85 -290 -65 -245
rect 670 -290 690 -245
rect 770 -290 790 5
rect 851 -61 871 83
rect 894 12 906 84
rect 928 12 937 84
rect 894 6 937 12
rect 959 86 1046 97
rect 1315 95 1337 133
rect 1575 150 1615 160
rect 1575 130 1585 150
rect 1605 130 1615 150
rect 1575 120 1615 130
rect 1790 150 1830 160
rect 1790 130 1800 150
rect 1820 130 1830 150
rect 1790 120 1830 130
rect 1953 144 1992 156
rect 1953 124 1963 144
rect 1983 124 1992 144
rect 1953 114 1992 124
rect 2070 134 2199 154
rect 2070 95 2089 134
rect 959 15 968 86
rect 989 74 1046 86
rect 989 15 1002 74
rect 959 6 1002 15
rect 895 -61 935 -60
rect 851 -70 935 -61
rect 851 -84 905 -70
rect 852 -86 905 -84
rect -250 -300 -210 -290
rect -250 -370 -240 -300
rect -220 -370 -210 -300
rect -250 -380 -210 -370
rect -170 -300 -130 -290
rect -170 -370 -160 -300
rect -140 -370 -130 -300
rect -170 -380 -130 -370
rect -105 -300 0 -290
rect -105 -370 -95 -300
rect -75 -370 -30 -300
rect -10 -370 0 -300
rect -105 -380 0 -370
rect 25 -300 65 -290
rect 25 -370 35 -300
rect 55 -370 65 -300
rect 25 -380 65 -370
rect 150 -300 190 -290
rect 150 -370 160 -300
rect 180 -370 190 -300
rect 150 -380 190 -370
rect 215 -300 255 -290
rect 215 -370 225 -300
rect 245 -370 255 -300
rect 215 -380 255 -370
rect 280 -300 325 -290
rect 280 -370 290 -300
rect 315 -370 325 -300
rect 280 -380 325 -370
rect 350 -300 390 -290
rect 350 -370 360 -300
rect 380 -370 390 -300
rect 350 -380 390 -370
rect 415 -300 455 -290
rect 415 -370 425 -300
rect 445 -370 455 -300
rect 415 -380 455 -370
rect 540 -300 580 -290
rect 540 -370 550 -300
rect 570 -370 580 -300
rect 540 -380 580 -370
rect 605 -300 710 -290
rect 605 -370 615 -300
rect 635 -370 680 -300
rect 700 -370 710 -300
rect 605 -380 710 -370
rect 735 -300 790 -290
rect 735 -370 745 -300
rect 765 -310 790 -300
rect 895 -140 905 -86
rect 925 -140 935 -70
rect 895 -225 935 -140
rect 960 -70 1000 -60
rect 960 -140 970 -70
rect 990 -140 1000 -70
rect 960 -150 1000 -140
rect 895 -295 905 -225
rect 925 -295 935 -225
rect 895 -305 935 -295
rect 959 -225 1000 -216
rect 959 -295 969 -225
rect 990 -295 1000 -225
rect 959 -306 1000 -295
rect 765 -370 775 -310
rect 1025 -344 1046 74
rect 1155 85 1195 95
rect 1155 15 1165 85
rect 1185 15 1195 85
rect 1250 85 1290 95
rect 1250 25 1260 85
rect 1155 5 1195 15
rect 1215 15 1260 25
rect 1280 15 1290 85
rect 1215 5 1290 15
rect 1315 85 1420 95
rect 1315 15 1325 85
rect 1345 15 1390 85
rect 1410 15 1420 85
rect 1315 5 1420 15
rect 1445 85 1485 95
rect 1445 15 1455 85
rect 1475 15 1485 85
rect 1445 5 1485 15
rect 1575 85 1615 95
rect 1575 15 1585 85
rect 1605 15 1615 85
rect 1575 5 1615 15
rect 1640 85 1680 95
rect 1640 15 1650 85
rect 1670 15 1680 85
rect 1640 5 1680 15
rect 1725 85 1765 95
rect 1725 15 1735 85
rect 1755 15 1765 85
rect 1725 5 1765 15
rect 1790 85 1830 95
rect 1790 15 1800 85
rect 1820 15 1830 85
rect 1790 5 1830 15
rect 1920 85 1960 95
rect 1920 15 1930 85
rect 1950 15 1960 85
rect 1920 5 1960 15
rect 1985 85 2090 95
rect 1985 15 1995 85
rect 2015 15 2060 85
rect 2080 15 2090 85
rect 1985 5 2090 15
rect 2115 85 2155 95
rect 2115 15 2125 85
rect 2145 25 2155 85
rect 2145 15 2190 25
rect 2115 5 2190 15
rect 1215 -255 1235 5
rect 1315 -15 1335 5
rect 1255 -35 1335 -15
rect 2070 -15 2090 5
rect 2070 -35 2150 -15
rect 1255 -205 1275 -35
rect 1485 -47 1920 -40
rect 1485 -66 1493 -47
rect 1512 -48 1920 -47
rect 1512 -60 1893 -48
rect 1512 -66 1520 -60
rect 1485 -75 1520 -66
rect 1590 -95 1610 -60
rect 1795 -95 1815 -60
rect 1885 -67 1893 -60
rect 1912 -67 1920 -48
rect 1885 -75 1920 -67
rect 1295 -105 1335 -95
rect 1295 -175 1305 -105
rect 1325 -175 1335 -105
rect 1295 -185 1335 -175
rect 1360 -105 1400 -95
rect 1360 -175 1370 -105
rect 1390 -175 1400 -105
rect 1360 -185 1400 -175
rect 1440 -105 1480 -95
rect 1440 -175 1450 -105
rect 1470 -175 1480 -105
rect 1440 -185 1480 -175
rect 1505 -105 1545 -95
rect 1505 -175 1515 -105
rect 1535 -175 1545 -105
rect 1505 -185 1545 -175
rect 1570 -105 1610 -95
rect 1570 -175 1580 -105
rect 1600 -175 1610 -105
rect 1570 -185 1610 -175
rect 1650 -105 1690 -95
rect 1650 -175 1660 -105
rect 1680 -175 1690 -105
rect 1650 -185 1690 -175
rect 1715 -105 1755 -95
rect 1715 -175 1725 -105
rect 1745 -175 1755 -105
rect 1715 -185 1755 -175
rect 1795 -105 1835 -95
rect 1795 -175 1805 -105
rect 1825 -175 1835 -105
rect 1795 -185 1835 -175
rect 1860 -105 1900 -95
rect 1860 -175 1870 -105
rect 1890 -175 1900 -105
rect 1860 -185 1900 -175
rect 1925 -105 1965 -95
rect 1925 -175 1935 -105
rect 1955 -175 1965 -105
rect 1925 -185 1965 -175
rect 2005 -105 2045 -95
rect 2005 -175 2015 -105
rect 2035 -175 2045 -105
rect 2005 -185 2045 -175
rect 2070 -105 2110 -95
rect 2070 -175 2080 -105
rect 2100 -175 2110 -105
rect 2070 -185 2110 -175
rect 1380 -205 1400 -185
rect 1735 -205 1755 -185
rect 2005 -205 2025 -185
rect 2130 -205 2150 -35
rect 1255 -215 1355 -205
rect 1255 -225 1325 -215
rect 1315 -235 1325 -225
rect 1345 -235 1355 -215
rect 1380 -225 2025 -205
rect 2050 -215 2150 -205
rect 1315 -245 1355 -235
rect 2050 -235 2060 -215
rect 2080 -225 2150 -215
rect 2080 -235 2090 -225
rect 2050 -245 2090 -235
rect 1215 -275 1250 -255
rect 1230 -290 1250 -275
rect 1315 -290 1335 -245
rect 2070 -290 2090 -245
rect 2170 -290 2190 5
rect 972 -345 1046 -344
rect 735 -380 775 -370
rect 894 -355 937 -345
rect -77 -407 -41 -398
rect -77 -427 -69 -407
rect -50 -417 -41 -407
rect 568 -407 604 -399
rect -50 -427 -38 -417
rect -77 -434 -38 -427
rect 568 -427 577 -407
rect 596 -427 604 -407
rect 568 -434 604 -427
rect -55 -435 604 -434
rect 894 -427 904 -355
rect 927 -427 937 -355
rect 894 -435 937 -427
rect 958 -356 1046 -345
rect 958 -427 967 -356
rect 988 -367 1046 -356
rect 1150 -300 1190 -290
rect 988 -427 1001 -367
rect 1150 -370 1160 -300
rect 1180 -370 1190 -300
rect 1150 -380 1190 -370
rect 1230 -300 1270 -290
rect 1230 -370 1240 -300
rect 1260 -370 1270 -300
rect 1230 -380 1270 -370
rect 1295 -300 1400 -290
rect 1295 -370 1305 -300
rect 1325 -370 1370 -300
rect 1390 -370 1400 -300
rect 1295 -380 1400 -370
rect 1425 -300 1465 -290
rect 1425 -370 1435 -300
rect 1455 -370 1465 -300
rect 1425 -380 1465 -370
rect 1550 -300 1590 -290
rect 1550 -370 1560 -300
rect 1580 -370 1590 -300
rect 1550 -380 1590 -370
rect 1615 -300 1655 -290
rect 1615 -370 1625 -300
rect 1645 -370 1655 -300
rect 1615 -380 1655 -370
rect 1680 -300 1725 -290
rect 1680 -370 1690 -300
rect 1715 -370 1725 -300
rect 1680 -380 1725 -370
rect 1750 -300 1790 -290
rect 1750 -370 1760 -300
rect 1780 -370 1790 -300
rect 1750 -380 1790 -370
rect 1815 -300 1855 -290
rect 1815 -370 1825 -300
rect 1845 -370 1855 -300
rect 1815 -380 1855 -370
rect 1940 -300 1980 -290
rect 1940 -370 1950 -300
rect 1970 -370 1980 -300
rect 1940 -380 1980 -370
rect 2005 -300 2110 -290
rect 2005 -370 2015 -300
rect 2035 -370 2080 -300
rect 2100 -370 2110 -300
rect 2005 -380 2110 -370
rect 2135 -300 2190 -290
rect 2135 -370 2145 -300
rect 2165 -310 2190 -300
rect 2165 -370 2175 -310
rect 2135 -380 2175 -370
rect 958 -435 1001 -427
rect 1323 -407 1359 -398
rect 1323 -427 1331 -407
rect 1350 -417 1359 -407
rect 1968 -407 2004 -399
rect 1350 -427 1362 -417
rect 1323 -434 1362 -427
rect 1968 -427 1977 -407
rect 1996 -427 2004 -407
rect 1968 -434 2004 -427
rect 1345 -435 2004 -434
rect -55 -453 586 -435
rect 1345 -453 1986 -435
rect -137 -463 -99 -455
rect -137 -485 -128 -463
rect -107 -473 -99 -463
rect 701 -464 740 -455
rect 701 -473 710 -464
rect -107 -485 710 -473
rect -137 -486 710 -485
rect 731 -486 740 -464
rect -137 -494 740 -486
rect 1263 -463 1301 -455
rect 1263 -485 1272 -463
rect 1293 -473 1301 -463
rect 2101 -464 2140 -455
rect 2101 -473 2110 -464
rect 1293 -485 2110 -473
rect 1263 -486 2110 -485
rect 2131 -486 2140 -464
rect 1263 -494 2140 -486
<< viali >>
rect -179 180 -156 205
rect 1221 180 1244 205
rect 185 130 205 150
rect 400 130 420 150
rect 563 124 583 144
rect -235 15 -215 85
rect 55 15 75 85
rect 185 15 205 85
rect 400 15 420 85
rect 530 15 550 85
rect -95 -175 -75 -105
rect 50 -175 70 -105
rect 115 -175 135 -105
rect 260 -175 280 -105
rect 470 -175 490 -105
rect 535 -175 555 -105
rect 680 -175 700 -105
rect 906 13 927 84
rect 927 13 928 84
rect 906 12 928 13
rect 1585 130 1605 150
rect 1800 130 1820 150
rect 1963 124 1983 144
rect -240 -370 -220 -300
rect 35 -370 55 -300
rect 160 -370 180 -300
rect 225 -370 245 -300
rect 360 -370 380 -300
rect 425 -370 445 -300
rect 550 -370 570 -300
rect 970 -140 990 -70
rect 969 -295 990 -225
rect 1165 15 1185 85
rect 1455 15 1475 85
rect 1585 15 1605 85
rect 1800 15 1820 85
rect 1930 15 1950 85
rect 1305 -175 1325 -105
rect 1450 -175 1470 -105
rect 1515 -175 1535 -105
rect 1660 -175 1680 -105
rect 1870 -175 1890 -105
rect 1935 -175 1955 -105
rect 2080 -175 2100 -105
rect 904 -356 927 -355
rect 904 -427 905 -356
rect 905 -427 926 -356
rect 926 -427 927 -356
rect 1160 -370 1180 -300
rect 1435 -370 1455 -300
rect 1560 -370 1580 -300
rect 1625 -370 1645 -300
rect 1760 -370 1780 -300
rect 1825 -370 1845 -300
rect 1950 -370 1970 -300
<< metal1 >>
rect -188 205 -146 214
rect -188 180 -179 205
rect -156 199 -146 205
rect 1212 205 1254 214
rect -7 199 576 200
rect -156 180 576 199
rect -188 177 576 180
rect 1212 180 1221 205
rect 1244 199 1254 205
rect 1393 199 1976 200
rect 1244 180 1976 199
rect 1212 177 1976 180
rect -188 175 30 177
rect -188 170 -146 175
rect 176 154 215 160
rect -165 150 215 154
rect -165 140 185 150
rect -245 85 -205 95
rect -245 15 -240 85
rect -210 15 -205 85
rect -245 5 -205 15
rect -250 -300 -210 -290
rect -250 -370 -245 -300
rect -215 -370 -210 -300
rect -250 -380 -210 -370
rect -165 -435 -135 140
rect 175 130 185 140
rect 205 130 215 150
rect 390 150 430 160
rect 559 156 575 177
rect 1212 175 1430 177
rect 1212 170 1254 175
rect 390 140 400 150
rect 175 120 215 130
rect 310 130 400 140
rect 420 130 430 150
rect 310 120 430 130
rect 552 144 592 156
rect 1576 154 1615 160
rect 552 124 563 144
rect 583 124 592 144
rect 45 85 85 95
rect 45 15 55 85
rect 75 15 85 85
rect 45 5 85 15
rect 175 90 215 95
rect 175 10 180 90
rect 210 10 215 90
rect 175 5 215 10
rect 45 -10 60 5
rect -15 -25 60 -10
rect -105 -105 -65 -95
rect -105 -175 -95 -105
rect -75 -175 -65 -105
rect -105 -185 -65 -175
rect -80 -400 -65 -185
rect -15 -290 0 -25
rect 40 -105 80 -95
rect 40 -175 50 -105
rect 70 -175 80 -105
rect 40 -185 80 -175
rect 105 -105 145 -95
rect 105 -175 115 -105
rect 135 -175 145 -105
rect 105 -185 145 -175
rect 250 -100 290 -95
rect 250 -180 255 -100
rect 285 -180 290 -100
rect 250 -185 290 -180
rect 65 -245 80 -185
rect 65 -260 230 -245
rect 215 -290 230 -260
rect -15 -300 65 -290
rect -15 -305 35 -300
rect 25 -370 35 -305
rect 55 -370 65 -300
rect 25 -380 65 -370
rect 150 -295 190 -290
rect 150 -375 155 -295
rect 185 -375 190 -295
rect 150 -380 190 -375
rect 215 -300 255 -290
rect 215 -370 225 -300
rect 245 -370 255 -300
rect 215 -380 255 -370
rect 310 -400 335 120
rect 552 113 592 124
rect 1235 150 1615 154
rect 1235 140 1585 150
rect 390 90 430 95
rect 390 10 395 90
rect 425 10 430 90
rect 390 5 430 10
rect 520 85 560 95
rect 520 15 530 85
rect 550 15 560 85
rect 520 5 560 15
rect 545 -10 560 5
rect 894 84 937 97
rect 894 12 906 84
rect 928 12 937 84
rect 545 -25 620 -10
rect 460 -105 500 -95
rect 460 -175 470 -105
rect 490 -175 500 -105
rect 460 -185 500 -175
rect 525 -105 565 -95
rect 525 -175 535 -105
rect 555 -175 565 -105
rect 525 -185 565 -175
rect 525 -250 540 -185
rect 375 -265 540 -250
rect 375 -290 390 -265
rect 605 -290 620 -25
rect 350 -300 390 -290
rect 350 -370 360 -300
rect 380 -370 390 -300
rect 350 -380 390 -370
rect 415 -295 455 -290
rect 415 -375 420 -295
rect 450 -375 455 -295
rect 415 -380 455 -375
rect 540 -300 620 -290
rect 540 -370 550 -300
rect 570 -305 620 -300
rect 670 -105 710 -95
rect 670 -175 680 -105
rect 700 -175 710 -105
rect 670 -185 710 -175
rect 570 -370 580 -305
rect 540 -380 580 -370
rect -80 -420 335 -400
rect 670 -435 690 -185
rect 894 -355 937 12
rect 1155 85 1195 95
rect 1155 15 1160 85
rect 1190 15 1195 85
rect 1155 5 1195 15
rect 960 -70 1000 -60
rect 960 -140 965 -70
rect 995 -140 1000 -70
rect 960 -150 1000 -140
rect 958 -224 1001 -216
rect 958 -295 964 -224
rect 995 -295 1001 -224
rect 958 -306 1001 -295
rect 1150 -300 1190 -290
rect 894 -427 904 -355
rect 927 -427 937 -355
rect 1150 -370 1155 -300
rect 1185 -370 1190 -300
rect 1150 -380 1190 -370
rect 894 -435 937 -427
rect 1235 -435 1265 140
rect 1575 130 1585 140
rect 1605 130 1615 150
rect 1790 150 1830 160
rect 1959 156 1975 177
rect 1790 140 1800 150
rect 1575 120 1615 130
rect 1710 130 1800 140
rect 1820 130 1830 150
rect 1710 120 1830 130
rect 1952 144 1992 156
rect 1952 124 1963 144
rect 1983 124 1992 144
rect 1445 85 1485 95
rect 1445 15 1455 85
rect 1475 15 1485 85
rect 1445 5 1485 15
rect 1575 90 1615 95
rect 1575 10 1580 90
rect 1610 10 1615 90
rect 1575 5 1615 10
rect 1445 -10 1460 5
rect 1385 -25 1460 -10
rect 1295 -105 1335 -95
rect 1295 -175 1305 -105
rect 1325 -175 1335 -105
rect 1295 -185 1335 -175
rect 1320 -400 1335 -185
rect 1385 -290 1400 -25
rect 1440 -105 1480 -95
rect 1440 -175 1450 -105
rect 1470 -175 1480 -105
rect 1440 -185 1480 -175
rect 1505 -105 1545 -95
rect 1505 -175 1515 -105
rect 1535 -175 1545 -105
rect 1505 -185 1545 -175
rect 1650 -100 1690 -95
rect 1650 -180 1655 -100
rect 1685 -180 1690 -100
rect 1650 -185 1690 -180
rect 1465 -245 1480 -185
rect 1465 -260 1630 -245
rect 1615 -290 1630 -260
rect 1385 -300 1465 -290
rect 1385 -305 1435 -300
rect 1425 -370 1435 -305
rect 1455 -370 1465 -300
rect 1425 -380 1465 -370
rect 1550 -295 1590 -290
rect 1550 -375 1555 -295
rect 1585 -375 1590 -295
rect 1550 -380 1590 -375
rect 1615 -300 1655 -290
rect 1615 -370 1625 -300
rect 1645 -370 1655 -300
rect 1615 -380 1655 -370
rect 1710 -400 1735 120
rect 1952 113 1992 124
rect 1790 90 1830 95
rect 1790 10 1795 90
rect 1825 10 1830 90
rect 1790 5 1830 10
rect 1920 85 1960 95
rect 1920 15 1930 85
rect 1950 15 1960 85
rect 1920 5 1960 15
rect 1945 -10 1960 5
rect 1945 -25 2020 -10
rect 1860 -105 1900 -95
rect 1860 -175 1870 -105
rect 1890 -175 1900 -105
rect 1860 -185 1900 -175
rect 1925 -105 1965 -95
rect 1925 -175 1935 -105
rect 1955 -175 1965 -105
rect 1925 -185 1965 -175
rect 1925 -250 1940 -185
rect 1775 -265 1940 -250
rect 1775 -290 1790 -265
rect 2005 -290 2020 -25
rect 1750 -300 1790 -290
rect 1750 -370 1760 -300
rect 1780 -370 1790 -300
rect 1750 -380 1790 -370
rect 1815 -295 1855 -290
rect 1815 -375 1820 -295
rect 1850 -375 1855 -295
rect 1815 -380 1855 -375
rect 1940 -300 2020 -290
rect 1940 -370 1950 -300
rect 1970 -305 2020 -300
rect 2070 -105 2110 -95
rect 2070 -175 2080 -105
rect 2100 -175 2110 -105
rect 2070 -185 2110 -175
rect 1970 -370 1980 -305
rect 1940 -380 1980 -370
rect 1320 -420 1735 -400
rect 2070 -435 2090 -185
rect -165 -455 690 -435
rect 1235 -455 2090 -435
<< via1 >>
rect -240 15 -235 85
rect -235 15 -215 85
rect -215 15 -210 85
rect -245 -370 -240 -300
rect -240 -370 -220 -300
rect -220 -370 -215 -300
rect 180 85 210 90
rect 180 15 185 85
rect 185 15 205 85
rect 205 15 210 85
rect 180 10 210 15
rect 255 -105 285 -100
rect 255 -175 260 -105
rect 260 -175 280 -105
rect 280 -175 285 -105
rect 255 -180 285 -175
rect 155 -300 185 -295
rect 155 -370 160 -300
rect 160 -370 180 -300
rect 180 -370 185 -300
rect 155 -375 185 -370
rect 395 85 425 90
rect 395 15 400 85
rect 400 15 420 85
rect 420 15 425 85
rect 395 10 425 15
rect 420 -300 450 -295
rect 420 -370 425 -300
rect 425 -370 445 -300
rect 445 -370 450 -300
rect 420 -375 450 -370
rect 1160 15 1165 85
rect 1165 15 1185 85
rect 1185 15 1190 85
rect 965 -140 970 -70
rect 970 -140 990 -70
rect 990 -140 995 -70
rect 964 -225 995 -224
rect 964 -295 969 -225
rect 969 -295 990 -225
rect 990 -295 995 -225
rect 1155 -370 1160 -300
rect 1160 -370 1180 -300
rect 1180 -370 1185 -300
rect 1580 85 1610 90
rect 1580 15 1585 85
rect 1585 15 1605 85
rect 1605 15 1610 85
rect 1580 10 1610 15
rect 1655 -105 1685 -100
rect 1655 -175 1660 -105
rect 1660 -175 1680 -105
rect 1680 -175 1685 -105
rect 1655 -180 1685 -175
rect 1555 -300 1585 -295
rect 1555 -370 1560 -300
rect 1560 -370 1580 -300
rect 1580 -370 1585 -300
rect 1555 -375 1585 -370
rect 1795 85 1825 90
rect 1795 15 1800 85
rect 1800 15 1820 85
rect 1820 15 1825 85
rect 1795 10 1825 15
rect 1820 -300 1850 -295
rect 1820 -370 1825 -300
rect 1825 -370 1845 -300
rect 1845 -370 1850 -300
rect 1820 -375 1850 -370
<< metal2 >>
rect -274 100 -188 101
rect 697 100 776 101
rect 2073 100 2201 101
rect -274 90 776 100
rect 1145 94 2201 100
rect -274 85 180 90
rect -274 15 -240 85
rect -210 15 180 85
rect -274 10 180 15
rect 210 10 395 90
rect 425 10 776 90
rect -274 0 776 10
rect 697 -45 776 0
rect 1141 90 2201 94
rect 1141 85 1580 90
rect 1141 15 1160 85
rect 1190 15 1580 85
rect 1141 10 1580 15
rect 1610 10 1795 90
rect 1825 10 2201 90
rect 1141 1 2201 10
rect 1141 0 2160 1
rect 1141 -45 1220 0
rect 697 -70 1220 -45
rect 250 -100 290 -95
rect 250 -180 255 -100
rect 285 -180 290 -100
rect 697 -140 965 -70
rect 995 -140 1220 -70
rect 697 -151 1220 -140
rect 1650 -100 1690 -95
rect 697 -152 776 -151
rect 955 -155 1005 -151
rect -273 -290 -107 -289
rect 250 -290 290 -180
rect 1650 -180 1655 -100
rect 1685 -180 1690 -100
rect 737 -224 1192 -207
rect 737 -290 964 -224
rect -273 -295 964 -290
rect 995 -290 1192 -224
rect 1650 -290 1690 -180
rect 995 -295 2201 -290
rect -273 -300 155 -295
rect -273 -370 -245 -300
rect -215 -370 155 -300
rect -273 -375 155 -370
rect 185 -375 420 -295
rect 450 -300 1555 -295
rect 450 -313 1155 -300
rect 450 -375 775 -313
rect -273 -380 775 -375
rect 1150 -370 1155 -313
rect 1185 -370 1555 -300
rect 1150 -375 1555 -370
rect 1585 -375 1820 -295
rect 1850 -375 2201 -295
rect 1150 -380 2201 -375
rect -263 -381 -107 -380
rect 2089 -382 2201 -380
<< labels >>
rlabel poly 300 145 300 145 5 Vb
port 1 s
rlabel poly 1700 145 1700 145 5 Vb
port 1 s
<< end >>
