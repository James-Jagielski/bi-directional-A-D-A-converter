magic
tech sky130A
timestamp 1702643716
<< nwell >>
rect 65 110 2070 250
rect 955 -20 1160 110
<< nmos >>
rect 135 -80 150 20
rect 200 -80 215 20
rect 410 -80 425 20
rect 475 -80 490 20
rect 540 -80 555 20
rect 605 -80 620 20
rect 815 -80 830 20
rect 1025 -155 1040 -55
rect 1305 -80 1320 20
rect 1515 -80 1530 20
rect 1580 -80 1595 20
rect 1645 -80 1660 20
rect 1710 -80 1725 20
rect 1920 -80 1935 20
rect 1985 -80 2000 20
rect 135 -275 150 -175
rect 200 -275 215 -175
rect 265 -275 280 -175
rect 410 -275 425 -175
rect 475 -275 490 -175
rect 540 -275 555 -175
rect 605 -275 620 -175
rect 750 -275 765 -175
rect 815 -275 830 -175
rect 880 -275 895 -175
rect 1025 -285 1040 -185
rect 1240 -275 1255 -175
rect 1305 -275 1320 -175
rect 1370 -275 1385 -175
rect 1515 -275 1530 -175
rect 1580 -275 1595 -175
rect 1645 -275 1660 -175
rect 1710 -275 1725 -175
rect 1855 -275 1870 -175
rect 1920 -275 1935 -175
rect 1985 -275 2000 -175
<< pmos >>
rect 135 130 150 230
rect 200 130 215 230
rect 265 130 280 230
rect 330 130 345 230
rect 370 130 385 230
rect 435 130 450 230
rect 580 130 595 230
rect 645 130 660 230
rect 685 130 700 230
rect 750 130 765 230
rect 815 130 830 230
rect 880 130 895 230
rect 1065 130 1080 230
rect 1240 130 1255 230
rect 1305 130 1320 230
rect 1370 130 1385 230
rect 1435 130 1450 230
rect 1475 130 1490 230
rect 1540 130 1555 230
rect 1685 130 1700 230
rect 1750 130 1765 230
rect 1790 130 1805 230
rect 1855 130 1870 230
rect 1920 130 1935 230
rect 1985 130 2000 230
rect 1025 0 1040 100
<< ndiff >>
rect 85 5 135 20
rect 85 -65 100 5
rect 120 -65 135 5
rect 85 -80 135 -65
rect 150 5 200 20
rect 150 -65 165 5
rect 185 -65 200 5
rect 150 -80 200 -65
rect 215 5 265 20
rect 215 -65 230 5
rect 250 -65 265 5
rect 215 -80 265 -65
rect 360 5 410 20
rect 360 -65 375 5
rect 395 -65 410 5
rect 360 -80 410 -65
rect 425 5 475 20
rect 425 -65 440 5
rect 460 -65 475 5
rect 425 -80 475 -65
rect 490 5 540 20
rect 490 -65 505 5
rect 525 -65 540 5
rect 490 -80 540 -65
rect 555 5 605 20
rect 555 -65 570 5
rect 590 -65 605 5
rect 555 -80 605 -65
rect 620 5 670 20
rect 620 -65 635 5
rect 655 -65 670 5
rect 620 -80 670 -65
rect 765 5 815 20
rect 765 -65 780 5
rect 800 -65 815 5
rect 765 -80 815 -65
rect 830 5 880 20
rect 830 -65 845 5
rect 865 -65 880 5
rect 1255 5 1305 20
rect 830 -80 880 -65
rect 975 -70 1025 -55
rect 975 -140 990 -70
rect 1010 -140 1025 -70
rect 975 -155 1025 -140
rect 1040 -70 1090 -55
rect 1040 -140 1055 -70
rect 1075 -140 1090 -70
rect 1255 -65 1270 5
rect 1290 -65 1305 5
rect 1255 -80 1305 -65
rect 1320 5 1370 20
rect 1320 -65 1335 5
rect 1355 -65 1370 5
rect 1320 -80 1370 -65
rect 1465 5 1515 20
rect 1465 -65 1480 5
rect 1500 -65 1515 5
rect 1465 -80 1515 -65
rect 1530 5 1580 20
rect 1530 -65 1545 5
rect 1565 -65 1580 5
rect 1530 -80 1580 -65
rect 1595 5 1645 20
rect 1595 -65 1610 5
rect 1630 -65 1645 5
rect 1595 -80 1645 -65
rect 1660 5 1710 20
rect 1660 -65 1675 5
rect 1695 -65 1710 5
rect 1660 -80 1710 -65
rect 1725 5 1775 20
rect 1725 -65 1740 5
rect 1760 -65 1775 5
rect 1725 -80 1775 -65
rect 1870 5 1920 20
rect 1870 -65 1885 5
rect 1905 -65 1920 5
rect 1870 -80 1920 -65
rect 1935 5 1985 20
rect 1935 -65 1950 5
rect 1970 -65 1985 5
rect 1935 -80 1985 -65
rect 2000 5 2050 20
rect 2000 -65 2015 5
rect 2035 -65 2050 5
rect 2000 -80 2050 -65
rect 1040 -155 1090 -140
rect 85 -190 135 -175
rect 85 -260 100 -190
rect 120 -260 135 -190
rect 85 -275 135 -260
rect 150 -190 200 -175
rect 150 -260 165 -190
rect 185 -260 200 -190
rect 150 -275 200 -260
rect 215 -190 265 -175
rect 215 -260 230 -190
rect 250 -260 265 -190
rect 215 -275 265 -260
rect 280 -190 330 -175
rect 280 -260 295 -190
rect 315 -260 330 -190
rect 280 -275 330 -260
rect 360 -190 410 -175
rect 360 -260 375 -190
rect 395 -260 410 -190
rect 360 -275 410 -260
rect 425 -190 475 -175
rect 425 -260 440 -190
rect 460 -260 475 -190
rect 425 -275 475 -260
rect 490 -190 540 -175
rect 490 -260 505 -190
rect 525 -260 540 -190
rect 490 -275 540 -260
rect 555 -190 605 -175
rect 555 -260 570 -190
rect 590 -260 605 -190
rect 555 -275 605 -260
rect 620 -190 670 -175
rect 620 -260 635 -190
rect 655 -260 670 -190
rect 620 -275 670 -260
rect 700 -190 750 -175
rect 700 -260 715 -190
rect 735 -260 750 -190
rect 700 -275 750 -260
rect 765 -190 815 -175
rect 765 -260 780 -190
rect 800 -260 815 -190
rect 765 -275 815 -260
rect 830 -190 880 -175
rect 830 -260 845 -190
rect 865 -260 880 -190
rect 830 -275 880 -260
rect 895 -190 945 -175
rect 895 -260 910 -190
rect 930 -260 945 -190
rect 895 -275 945 -260
rect 975 -200 1025 -185
rect 975 -270 990 -200
rect 1010 -270 1025 -200
rect 975 -285 1025 -270
rect 1040 -200 1090 -185
rect 1040 -270 1055 -200
rect 1075 -270 1090 -200
rect 1040 -285 1090 -270
rect 1190 -190 1240 -175
rect 1190 -260 1205 -190
rect 1225 -260 1240 -190
rect 1190 -275 1240 -260
rect 1255 -190 1305 -175
rect 1255 -260 1270 -190
rect 1290 -260 1305 -190
rect 1255 -275 1305 -260
rect 1320 -190 1370 -175
rect 1320 -260 1335 -190
rect 1355 -260 1370 -190
rect 1320 -275 1370 -260
rect 1385 -190 1435 -175
rect 1385 -260 1400 -190
rect 1420 -260 1435 -190
rect 1385 -275 1435 -260
rect 1465 -190 1515 -175
rect 1465 -260 1480 -190
rect 1500 -260 1515 -190
rect 1465 -275 1515 -260
rect 1530 -190 1580 -175
rect 1530 -260 1545 -190
rect 1565 -260 1580 -190
rect 1530 -275 1580 -260
rect 1595 -190 1645 -175
rect 1595 -260 1610 -190
rect 1630 -260 1645 -190
rect 1595 -275 1645 -260
rect 1660 -190 1710 -175
rect 1660 -260 1675 -190
rect 1695 -260 1710 -190
rect 1660 -275 1710 -260
rect 1725 -190 1775 -175
rect 1725 -260 1740 -190
rect 1760 -260 1775 -190
rect 1725 -275 1775 -260
rect 1805 -190 1855 -175
rect 1805 -260 1820 -190
rect 1840 -260 1855 -190
rect 1805 -275 1855 -260
rect 1870 -190 1920 -175
rect 1870 -260 1885 -190
rect 1905 -260 1920 -190
rect 1870 -275 1920 -260
rect 1935 -190 1985 -175
rect 1935 -260 1950 -190
rect 1970 -260 1985 -190
rect 1935 -275 1985 -260
rect 2000 -190 2050 -175
rect 2000 -260 2015 -190
rect 2035 -260 2050 -190
rect 2000 -275 2050 -260
<< pdiff >>
rect 85 215 135 230
rect 85 145 100 215
rect 120 145 135 215
rect 85 130 135 145
rect 150 215 200 230
rect 150 145 165 215
rect 185 145 200 215
rect 150 130 200 145
rect 215 215 265 230
rect 215 145 230 215
rect 250 145 265 215
rect 215 130 265 145
rect 280 215 330 230
rect 280 145 295 215
rect 315 145 330 215
rect 280 130 330 145
rect 345 130 370 230
rect 385 215 435 230
rect 385 145 400 215
rect 420 145 435 215
rect 385 130 435 145
rect 450 215 500 230
rect 450 145 465 215
rect 485 145 500 215
rect 450 130 500 145
rect 530 215 580 230
rect 530 145 545 215
rect 565 145 580 215
rect 530 130 580 145
rect 595 215 645 230
rect 595 145 610 215
rect 630 145 645 215
rect 595 130 645 145
rect 660 130 685 230
rect 700 215 750 230
rect 700 145 715 215
rect 735 145 750 215
rect 700 130 750 145
rect 765 215 815 230
rect 765 145 780 215
rect 800 145 815 215
rect 765 130 815 145
rect 830 215 880 230
rect 830 145 845 215
rect 865 145 880 215
rect 830 130 880 145
rect 895 215 945 230
rect 895 145 910 215
rect 930 145 945 215
rect 1015 215 1065 230
rect 895 130 945 145
rect 1015 145 1030 215
rect 1050 145 1065 215
rect 1015 130 1065 145
rect 1080 215 1130 230
rect 1080 145 1095 215
rect 1115 145 1130 215
rect 1080 130 1130 145
rect 1190 215 1240 230
rect 1190 145 1205 215
rect 1225 145 1240 215
rect 1190 130 1240 145
rect 1255 215 1305 230
rect 1255 145 1270 215
rect 1290 145 1305 215
rect 1255 130 1305 145
rect 1320 215 1370 230
rect 1320 145 1335 215
rect 1355 145 1370 215
rect 1320 130 1370 145
rect 1385 215 1435 230
rect 1385 145 1400 215
rect 1420 145 1435 215
rect 1385 130 1435 145
rect 1450 130 1475 230
rect 1490 215 1540 230
rect 1490 145 1505 215
rect 1525 145 1540 215
rect 1490 130 1540 145
rect 1555 215 1605 230
rect 1555 145 1570 215
rect 1590 145 1605 215
rect 1555 130 1605 145
rect 1635 215 1685 230
rect 1635 145 1650 215
rect 1670 145 1685 215
rect 1635 130 1685 145
rect 1700 215 1750 230
rect 1700 145 1715 215
rect 1735 145 1750 215
rect 1700 130 1750 145
rect 1765 130 1790 230
rect 1805 215 1855 230
rect 1805 145 1820 215
rect 1840 145 1855 215
rect 1805 130 1855 145
rect 1870 215 1920 230
rect 1870 145 1885 215
rect 1905 145 1920 215
rect 1870 130 1920 145
rect 1935 215 1985 230
rect 1935 145 1950 215
rect 1970 145 1985 215
rect 1935 130 1985 145
rect 2000 215 2050 230
rect 2000 145 2015 215
rect 2035 145 2050 215
rect 2000 130 2050 145
rect 975 85 1025 100
rect 975 15 990 85
rect 1010 15 1025 85
rect 975 0 1025 15
rect 1040 85 1090 100
rect 1040 15 1055 85
rect 1075 15 1090 85
rect 1040 0 1090 15
<< ndiffc >>
rect 100 -65 120 5
rect 165 -65 185 5
rect 230 -65 250 5
rect 375 -65 395 5
rect 440 -65 460 5
rect 505 -65 525 5
rect 570 -65 590 5
rect 635 -65 655 5
rect 780 -65 800 5
rect 845 -65 865 5
rect 990 -140 1010 -70
rect 1055 -140 1075 -70
rect 1270 -65 1290 5
rect 1335 -65 1355 5
rect 1480 -65 1500 5
rect 1545 -65 1565 5
rect 1610 -65 1630 5
rect 1675 -65 1695 5
rect 1740 -65 1760 5
rect 1885 -65 1905 5
rect 1950 -65 1970 5
rect 2015 -65 2035 5
rect 100 -260 120 -190
rect 165 -260 185 -190
rect 230 -260 250 -190
rect 295 -260 315 -190
rect 375 -260 395 -190
rect 440 -260 460 -190
rect 505 -260 525 -190
rect 570 -260 590 -190
rect 635 -260 655 -190
rect 715 -260 735 -190
rect 780 -260 800 -190
rect 845 -260 865 -190
rect 910 -260 930 -190
rect 990 -270 1010 -200
rect 1055 -270 1075 -200
rect 1205 -260 1225 -190
rect 1270 -260 1290 -190
rect 1335 -260 1355 -190
rect 1400 -260 1420 -190
rect 1480 -260 1500 -190
rect 1545 -260 1565 -190
rect 1610 -260 1630 -190
rect 1675 -260 1695 -190
rect 1740 -260 1760 -190
rect 1820 -260 1840 -190
rect 1885 -260 1905 -190
rect 1950 -260 1970 -190
rect 2015 -260 2035 -190
<< pdiffc >>
rect 100 145 120 215
rect 165 145 185 215
rect 230 145 250 215
rect 295 145 315 215
rect 400 145 420 215
rect 465 145 485 215
rect 545 145 565 215
rect 610 145 630 215
rect 715 145 735 215
rect 780 145 800 215
rect 845 145 865 215
rect 910 145 930 215
rect 1030 145 1050 215
rect 1095 145 1115 215
rect 1205 145 1225 215
rect 1270 145 1290 215
rect 1335 145 1355 215
rect 1400 145 1420 215
rect 1505 145 1525 215
rect 1570 145 1590 215
rect 1650 145 1670 215
rect 1715 145 1735 215
rect 1820 145 1840 215
rect 1885 145 1905 215
rect 1950 145 1970 215
rect 2015 145 2035 215
rect 990 15 1010 85
rect 1055 15 1075 85
<< psubdiff >>
rect 1090 -70 1140 -55
rect 1090 -140 1105 -70
rect 1125 -140 1140 -70
rect 1090 -155 1140 -140
<< nsubdiff >>
rect 1090 85 1140 100
rect 1090 15 1105 85
rect 1125 15 1140 85
rect 1090 0 1140 15
<< psubdiffcont >>
rect 1105 -140 1125 -70
<< nsubdiffcont >>
rect 1105 15 1125 85
<< poly >>
rect 775 390 895 405
rect 775 365 790 390
rect 135 350 790 365
rect 815 355 855 365
rect 135 230 150 350
rect 815 335 825 355
rect 845 335 855 355
rect 815 325 855 335
rect 200 315 790 325
rect 200 310 760 315
rect 200 230 215 310
rect 750 295 760 310
rect 780 295 790 315
rect 750 285 790 295
rect 265 275 305 285
rect 265 255 275 275
rect 295 255 305 275
rect 265 245 305 255
rect 330 275 725 285
rect 330 270 695 275
rect 265 230 280 245
rect 330 230 345 270
rect 685 255 695 270
rect 715 255 725 275
rect 685 245 725 255
rect 370 230 385 245
rect 435 230 450 245
rect 580 230 595 245
rect 645 230 660 245
rect 685 230 700 245
rect 750 230 765 285
rect 815 230 830 325
rect 880 300 895 390
rect 1240 350 2000 365
rect 1240 300 1255 350
rect 880 285 1255 300
rect 1280 315 1320 325
rect 1280 295 1290 315
rect 1310 295 1320 315
rect 1280 285 1320 295
rect 880 230 895 285
rect 985 245 1080 260
rect 985 220 1000 245
rect 1065 230 1080 245
rect 1240 230 1255 285
rect 1305 230 1320 285
rect 1370 315 1935 325
rect 1370 310 1905 315
rect 1370 230 1385 310
rect 1895 295 1905 310
rect 1925 295 1935 315
rect 1895 285 1935 295
rect 1410 275 1805 285
rect 1410 255 1420 275
rect 1440 270 1805 275
rect 1440 255 1450 270
rect 1410 245 1450 255
rect 1435 230 1450 245
rect 1475 230 1490 245
rect 1540 230 1555 245
rect 1685 230 1700 245
rect 1750 230 1765 245
rect 1790 230 1805 270
rect 1830 275 1870 285
rect 1830 255 1840 275
rect 1860 255 1870 275
rect 1830 245 1870 255
rect 1855 230 1870 245
rect 1920 230 1935 285
rect 1985 230 2000 350
rect 960 210 1000 220
rect 960 190 970 210
rect 990 190 1000 210
rect 960 180 1000 190
rect 135 115 150 130
rect 200 115 215 130
rect 265 115 280 130
rect 330 115 345 130
rect 370 115 385 130
rect 435 115 450 130
rect 370 105 450 115
rect 200 80 240 90
rect 135 65 175 75
rect 135 45 145 65
rect 165 45 175 65
rect 135 35 175 45
rect 200 60 210 80
rect 230 60 240 80
rect 370 85 380 105
rect 400 100 450 105
rect 580 115 595 130
rect 645 115 660 130
rect 685 115 700 130
rect 750 115 765 130
rect 815 115 830 130
rect 880 115 895 130
rect 1065 115 1080 130
rect 1240 115 1255 130
rect 1305 115 1320 130
rect 1370 115 1385 130
rect 1435 115 1450 130
rect 1475 115 1490 130
rect 1540 115 1555 130
rect 580 105 660 115
rect 580 100 630 105
rect 400 85 410 100
rect 370 75 410 85
rect 620 85 630 100
rect 650 85 660 105
rect 1025 100 1040 115
rect 1475 105 1555 115
rect 620 75 660 85
rect 200 50 240 60
rect 455 65 495 75
rect 135 20 150 35
rect 200 20 215 50
rect 455 45 465 65
rect 485 45 495 65
rect 455 35 495 45
rect 535 65 575 75
rect 535 45 545 65
rect 565 45 575 65
rect 535 35 575 45
rect 410 20 425 35
rect 475 20 490 35
rect 540 20 555 35
rect 605 20 620 35
rect 815 20 830 35
rect 1475 85 1485 105
rect 1505 100 1555 105
rect 1685 115 1700 130
rect 1750 115 1765 130
rect 1790 115 1805 130
rect 1855 115 1870 130
rect 1920 115 1935 130
rect 1985 115 2000 130
rect 1685 105 1765 115
rect 1685 100 1735 105
rect 1505 85 1515 100
rect 1475 75 1515 85
rect 1725 85 1735 100
rect 1755 85 1765 105
rect 1725 75 1765 85
rect 1560 65 1600 75
rect 1560 45 1570 65
rect 1590 45 1600 65
rect 1560 35 1600 45
rect 1640 65 1680 75
rect 1640 45 1650 65
rect 1670 45 1680 65
rect 1640 35 1680 45
rect 1895 65 1935 75
rect 1895 45 1905 65
rect 1925 45 1935 65
rect 1895 35 1935 45
rect 1960 65 2000 75
rect 1960 45 1970 65
rect 1990 45 2000 65
rect 1960 35 2000 45
rect 1305 20 1320 35
rect 1515 20 1530 35
rect 1580 20 1595 35
rect 1645 20 1660 35
rect 1710 20 1725 35
rect 1920 20 1935 35
rect 1985 20 2000 35
rect 1025 -55 1040 0
rect 135 -95 150 -80
rect 200 -95 215 -80
rect 410 -95 425 -80
rect 135 -105 175 -95
rect 135 -125 145 -105
rect 165 -125 175 -105
rect 135 -135 175 -125
rect 410 -105 450 -95
rect 410 -125 420 -105
rect 440 -125 450 -105
rect 410 -135 450 -125
rect 135 -175 150 -160
rect 200 -175 215 -160
rect 265 -175 280 -160
rect 410 -175 425 -160
rect 475 -175 490 -80
rect 540 -175 555 -80
rect 605 -95 620 -80
rect 815 -95 830 -80
rect 580 -105 620 -95
rect 580 -125 590 -105
rect 610 -125 620 -105
rect 580 -135 620 -125
rect 790 -105 830 -95
rect 790 -125 800 -105
rect 820 -125 830 -105
rect 790 -135 830 -125
rect 1305 -95 1320 -80
rect 1515 -95 1530 -80
rect 1305 -105 1345 -95
rect 1305 -125 1315 -105
rect 1335 -125 1345 -105
rect 1305 -135 1345 -125
rect 1515 -105 1555 -95
rect 1515 -125 1525 -105
rect 1545 -125 1555 -105
rect 1515 -135 1555 -125
rect 605 -175 620 -160
rect 750 -175 765 -160
rect 815 -175 830 -160
rect 880 -175 895 -160
rect 1025 -185 1040 -155
rect 1240 -175 1255 -160
rect 1305 -175 1320 -160
rect 1370 -175 1385 -160
rect 1515 -175 1530 -160
rect 1580 -175 1595 -80
rect 1645 -175 1660 -80
rect 1710 -95 1725 -80
rect 1920 -95 1935 -80
rect 1985 -95 2000 -80
rect 1685 -105 1725 -95
rect 1685 -125 1695 -105
rect 1715 -125 1725 -105
rect 1685 -135 1725 -125
rect 1960 -105 2000 -95
rect 1960 -125 1970 -105
rect 1990 -125 2000 -105
rect 1960 -135 2000 -125
rect 1710 -175 1725 -160
rect 1855 -175 1870 -160
rect 1920 -175 1935 -160
rect 1985 -175 2000 -160
rect 135 -395 150 -275
rect 200 -290 215 -275
rect 200 -300 240 -290
rect 200 -320 210 -300
rect 230 -320 240 -300
rect 200 -330 240 -320
rect 265 -355 280 -275
rect 410 -315 425 -275
rect 475 -290 490 -275
rect 540 -290 555 -275
rect 605 -290 620 -275
rect 750 -290 765 -275
rect 580 -300 620 -290
rect 580 -315 590 -300
rect 410 -320 590 -315
rect 610 -320 620 -300
rect 410 -330 620 -320
rect 715 -300 765 -290
rect 715 -320 725 -300
rect 745 -305 765 -300
rect 745 -320 755 -305
rect 715 -330 755 -320
rect 815 -330 830 -275
rect 780 -340 830 -330
rect 780 -355 790 -340
rect 265 -360 790 -355
rect 810 -345 830 -340
rect 810 -360 820 -345
rect 265 -370 820 -360
rect 880 -395 895 -275
rect 1025 -300 1040 -285
rect 1240 -395 1255 -275
rect 1305 -290 1320 -275
rect 1305 -300 1345 -290
rect 1305 -320 1315 -300
rect 1335 -320 1345 -300
rect 1305 -330 1345 -320
rect 1370 -330 1385 -275
rect 1515 -290 1530 -275
rect 1580 -290 1595 -275
rect 1645 -290 1660 -275
rect 1515 -300 1555 -290
rect 1515 -320 1525 -300
rect 1545 -315 1555 -300
rect 1710 -315 1725 -275
rect 1855 -290 1870 -275
rect 1545 -320 1725 -315
rect 1515 -330 1725 -320
rect 1830 -300 1870 -290
rect 1830 -320 1840 -300
rect 1860 -320 1870 -300
rect 1830 -330 1870 -320
rect 1370 -340 1410 -330
rect 1370 -360 1380 -340
rect 1400 -355 1410 -340
rect 1920 -355 1935 -275
rect 1400 -360 1935 -355
rect 1370 -370 1935 -360
rect 1985 -395 2000 -275
rect 135 -410 2000 -395
<< polycont >>
rect 825 335 845 355
rect 760 295 780 315
rect 275 255 295 275
rect 695 255 715 275
rect 1290 295 1310 315
rect 1905 295 1925 315
rect 1420 255 1440 275
rect 1840 255 1860 275
rect 970 190 990 210
rect 145 45 165 65
rect 210 60 230 80
rect 380 85 400 105
rect 630 85 650 105
rect 465 45 485 65
rect 545 45 565 65
rect 1485 85 1505 105
rect 1735 85 1755 105
rect 1570 45 1590 65
rect 1650 45 1670 65
rect 1905 45 1925 65
rect 1970 45 1990 65
rect 145 -125 165 -105
rect 420 -125 440 -105
rect 590 -125 610 -105
rect 800 -125 820 -105
rect 1315 -125 1335 -105
rect 1525 -125 1545 -105
rect 1695 -125 1715 -105
rect 1970 -125 1990 -105
rect 210 -320 230 -300
rect 590 -320 610 -300
rect 725 -320 745 -300
rect 790 -360 810 -340
rect 1315 -320 1335 -300
rect 1525 -320 1545 -300
rect 1840 -320 1860 -300
rect 1380 -360 1400 -340
<< locali >>
rect 640 355 1530 365
rect 640 345 825 355
rect 640 285 660 345
rect 815 335 825 345
rect 845 345 1530 355
rect 845 335 855 345
rect 815 325 855 335
rect 1510 325 1530 345
rect 750 315 790 325
rect 750 295 760 315
rect 780 305 790 315
rect 1280 315 1490 325
rect 1280 305 1290 315
rect 780 295 1290 305
rect 1310 305 1490 315
rect 1510 315 1935 325
rect 1510 305 1905 315
rect 1310 295 1320 305
rect 750 285 1320 295
rect 265 275 660 285
rect 265 255 275 275
rect 295 265 660 275
rect 685 275 725 285
rect 295 255 305 265
rect 265 245 305 255
rect 685 255 695 275
rect 715 265 725 275
rect 1410 275 1450 285
rect 1410 265 1420 275
rect 715 255 1420 265
rect 1440 255 1450 275
rect 685 245 1450 255
rect 1470 265 1490 305
rect 1895 295 1905 305
rect 1925 295 1935 315
rect 1895 285 1935 295
rect 1830 275 1870 285
rect 1830 265 1840 275
rect 1470 255 1840 265
rect 1860 255 1870 275
rect 1470 245 1870 255
rect 90 215 130 225
rect 90 155 100 215
rect 50 145 100 155
rect 120 145 130 215
rect 50 135 130 145
rect 155 215 260 225
rect 155 145 165 215
rect 185 145 230 215
rect 250 145 260 215
rect 155 135 260 145
rect 285 215 325 225
rect 285 145 295 215
rect 315 145 325 215
rect 50 -180 70 135
rect 155 75 175 135
rect 135 65 175 75
rect 135 45 145 65
rect 165 45 175 65
rect 200 60 210 90
rect 230 60 240 90
rect 200 50 240 60
rect 135 35 175 45
rect 90 5 130 15
rect 90 -65 100 5
rect 120 -65 130 5
rect 90 -75 130 -65
rect 155 5 195 15
rect 155 -65 165 5
rect 185 -65 195 5
rect 155 -75 195 -65
rect 220 5 260 15
rect 220 -65 230 5
rect 250 -65 260 5
rect 220 -75 260 -65
rect 285 -45 325 145
rect 390 215 430 225
rect 390 145 400 215
rect 420 145 430 215
rect 390 135 430 145
rect 455 215 495 225
rect 455 145 465 215
rect 485 145 495 215
rect 455 135 495 145
rect 535 215 575 225
rect 535 145 545 215
rect 565 145 575 215
rect 535 135 575 145
rect 600 215 640 225
rect 600 145 610 215
rect 630 145 640 215
rect 600 135 640 145
rect 705 215 745 225
rect 705 145 715 215
rect 735 145 745 215
rect 705 135 745 145
rect 770 215 875 225
rect 770 145 780 215
rect 800 145 845 215
rect 865 145 875 215
rect 770 135 875 145
rect 900 215 940 225
rect 900 145 910 215
rect 930 155 940 215
rect 960 210 1000 220
rect 960 190 970 210
rect 990 190 1000 210
rect 960 180 1000 190
rect 930 145 955 155
rect 900 135 955 145
rect 455 115 475 135
rect 370 105 475 115
rect 370 85 380 105
rect 400 95 475 105
rect 555 115 575 135
rect 555 105 660 115
rect 555 95 630 105
rect 400 85 410 95
rect 370 75 410 85
rect 620 85 630 95
rect 650 95 660 105
rect 650 85 695 95
rect 620 75 695 85
rect 455 70 495 75
rect 455 45 465 70
rect 485 45 495 70
rect 455 35 495 45
rect 535 70 575 75
rect 535 45 545 70
rect 565 45 575 70
rect 535 35 575 45
rect 675 60 695 75
rect 675 55 705 60
rect 675 35 680 55
rect 700 35 705 55
rect 675 30 705 35
rect 285 -65 295 -45
rect 315 -65 325 -45
rect 135 -105 175 -95
rect 135 -125 145 -105
rect 165 -125 175 -105
rect 135 -135 175 -125
rect 155 -180 175 -135
rect 50 -190 130 -180
rect 50 -200 100 -190
rect 90 -260 100 -200
rect 120 -260 130 -190
rect 90 -270 130 -260
rect 155 -190 260 -180
rect 155 -260 165 -190
rect 185 -260 230 -190
rect 250 -260 260 -190
rect 155 -270 260 -260
rect 285 -190 325 -65
rect 365 5 405 15
rect 365 -65 375 5
rect 395 -65 405 5
rect 365 -75 405 -65
rect 430 5 470 15
rect 430 -65 440 5
rect 460 -65 470 5
rect 430 -75 470 -65
rect 495 5 535 15
rect 495 -65 505 5
rect 525 -65 535 5
rect 365 -120 385 -75
rect 495 -95 535 -65
rect 560 5 600 15
rect 560 -65 570 5
rect 590 -65 600 5
rect 560 -75 600 -65
rect 625 5 665 15
rect 625 -65 635 5
rect 655 -65 665 5
rect 725 -35 745 135
rect 855 110 875 135
rect 855 100 915 110
rect 855 90 885 100
rect 875 80 885 90
rect 905 80 915 100
rect 875 70 915 80
rect 625 -75 665 -65
rect 345 -130 385 -120
rect 345 -150 355 -130
rect 375 -150 385 -130
rect 410 -105 620 -95
rect 410 -125 420 -105
rect 440 -115 590 -105
rect 440 -125 450 -115
rect 410 -135 450 -125
rect 580 -125 590 -115
rect 610 -125 620 -105
rect 580 -135 620 -125
rect 645 -120 665 -75
rect 705 -45 745 -35
rect 705 -65 715 -45
rect 735 -65 745 -45
rect 645 -130 685 -120
rect 345 -160 385 -150
rect 645 -150 655 -130
rect 675 -150 685 -130
rect 645 -160 685 -150
rect 285 -260 295 -190
rect 315 -260 325 -190
rect 285 -270 325 -260
rect 365 -190 405 -180
rect 365 -260 375 -190
rect 395 -260 405 -190
rect 365 -270 405 -260
rect 430 -190 470 -180
rect 430 -260 440 -190
rect 460 -260 470 -190
rect 430 -270 470 -260
rect 495 -190 535 -180
rect 495 -260 505 -190
rect 525 -260 535 -190
rect 495 -270 535 -260
rect 560 -190 600 -180
rect 560 -260 570 -190
rect 590 -260 600 -190
rect 560 -270 600 -260
rect 625 -190 665 -180
rect 625 -260 635 -190
rect 655 -260 665 -190
rect 625 -270 665 -260
rect 705 -190 745 -65
rect 770 5 810 15
rect 770 -65 780 5
rect 800 -65 810 5
rect 770 -75 810 -65
rect 835 5 875 15
rect 835 -65 845 5
rect 865 -65 875 5
rect 835 -75 875 -65
rect 895 -95 915 70
rect 790 -105 915 -95
rect 790 -125 800 -105
rect 820 -115 915 -105
rect 820 -125 830 -115
rect 790 -180 830 -125
rect 935 -180 955 135
rect 980 95 1000 180
rect 1020 215 1060 225
rect 1020 145 1030 215
rect 1050 145 1060 215
rect 1020 135 1060 145
rect 1085 215 1125 225
rect 1085 145 1095 215
rect 1115 155 1125 215
rect 1195 215 1235 225
rect 1115 145 1175 155
rect 1085 135 1175 145
rect 1195 145 1205 215
rect 1225 145 1235 215
rect 1195 135 1235 145
rect 1260 215 1365 225
rect 1260 145 1270 215
rect 1290 145 1335 215
rect 1355 145 1365 215
rect 1260 135 1365 145
rect 1390 215 1430 225
rect 1390 145 1400 215
rect 1420 145 1430 215
rect 1390 135 1430 145
rect 1495 215 1535 225
rect 1495 145 1505 215
rect 1525 145 1535 215
rect 1495 135 1535 145
rect 1560 215 1600 225
rect 1560 145 1570 215
rect 1590 145 1600 215
rect 1560 135 1600 145
rect 1640 215 1680 225
rect 1640 145 1650 215
rect 1670 145 1680 215
rect 1640 135 1680 145
rect 1705 215 1745 225
rect 1705 145 1715 215
rect 1735 145 1745 215
rect 1705 135 1745 145
rect 1810 215 1850 225
rect 1810 145 1820 215
rect 1840 145 1850 215
rect 1155 110 1175 135
rect 1260 110 1280 135
rect 980 85 1020 95
rect 980 15 990 85
rect 1010 15 1020 85
rect 980 -70 1020 15
rect 1045 85 1135 95
rect 1155 90 1280 110
rect 1045 15 1055 85
rect 1075 15 1105 85
rect 1125 15 1135 85
rect 1045 5 1135 15
rect 980 -140 990 -70
rect 1010 -140 1020 -70
rect 980 -150 1020 -140
rect 1045 -70 1135 -60
rect 1045 -140 1055 -70
rect 1075 -140 1105 -70
rect 1125 -140 1135 -70
rect 1220 -95 1240 90
rect 1260 5 1300 15
rect 1260 -65 1270 5
rect 1290 -65 1300 5
rect 1260 -75 1300 -65
rect 1325 5 1365 15
rect 1325 -65 1335 5
rect 1355 -65 1365 5
rect 1325 -75 1365 -65
rect 1390 -35 1410 135
rect 1560 115 1580 135
rect 1475 105 1580 115
rect 1475 95 1485 105
rect 1440 85 1485 95
rect 1505 95 1580 105
rect 1660 115 1680 135
rect 1660 105 1765 115
rect 1660 95 1735 105
rect 1505 85 1515 95
rect 1440 75 1515 85
rect 1725 85 1735 95
rect 1755 85 1765 105
rect 1725 75 1765 85
rect 1440 60 1460 75
rect 1430 55 1460 60
rect 1430 35 1435 55
rect 1455 35 1460 55
rect 1560 70 1600 75
rect 1560 45 1570 70
rect 1590 45 1600 70
rect 1560 35 1600 45
rect 1640 70 1680 75
rect 1640 45 1650 70
rect 1670 45 1680 70
rect 1640 35 1680 45
rect 1430 30 1460 35
rect 1470 5 1510 15
rect 1390 -45 1430 -35
rect 1390 -65 1400 -45
rect 1420 -65 1430 -45
rect 1045 -150 1135 -140
rect 1155 -105 1345 -95
rect 1155 -115 1315 -105
rect 705 -260 715 -190
rect 735 -260 745 -190
rect 705 -270 745 -260
rect 770 -190 875 -180
rect 770 -260 780 -190
rect 800 -260 845 -190
rect 865 -260 875 -190
rect 770 -270 875 -260
rect 900 -190 955 -180
rect 1155 -190 1175 -115
rect 1305 -125 1315 -115
rect 1335 -125 1345 -105
rect 1305 -180 1345 -125
rect 900 -260 910 -190
rect 930 -200 955 -190
rect 980 -200 1020 -190
rect 930 -260 940 -200
rect 900 -270 940 -260
rect 980 -270 990 -200
rect 1010 -270 1020 -200
rect 515 -290 535 -270
rect 980 -280 1020 -270
rect 1045 -200 1175 -190
rect 1045 -270 1055 -200
rect 1075 -210 1175 -200
rect 1195 -190 1235 -180
rect 1075 -270 1085 -210
rect 1195 -260 1205 -190
rect 1225 -260 1235 -190
rect 1195 -270 1235 -260
rect 1260 -190 1365 -180
rect 1260 -260 1270 -190
rect 1290 -260 1335 -190
rect 1355 -260 1365 -190
rect 1260 -270 1365 -260
rect 1390 -190 1430 -65
rect 1470 -65 1480 5
rect 1500 -65 1510 5
rect 1470 -75 1510 -65
rect 1535 5 1575 15
rect 1535 -65 1545 5
rect 1565 -65 1575 5
rect 1535 -75 1575 -65
rect 1600 5 1640 15
rect 1600 -65 1610 5
rect 1630 -65 1640 5
rect 1470 -120 1490 -75
rect 1600 -95 1640 -65
rect 1665 5 1705 15
rect 1665 -65 1675 5
rect 1695 -65 1705 5
rect 1665 -75 1705 -65
rect 1730 5 1770 15
rect 1730 -65 1740 5
rect 1760 -65 1770 5
rect 1730 -75 1770 -65
rect 1450 -130 1490 -120
rect 1450 -150 1460 -130
rect 1480 -150 1490 -130
rect 1515 -105 1725 -95
rect 1515 -125 1525 -105
rect 1545 -115 1695 -105
rect 1545 -125 1555 -115
rect 1515 -135 1555 -125
rect 1685 -125 1695 -115
rect 1715 -125 1725 -105
rect 1685 -135 1725 -125
rect 1750 -120 1770 -75
rect 1810 -45 1850 145
rect 1875 215 1980 225
rect 1875 145 1885 215
rect 1905 145 1950 215
rect 1970 145 1980 215
rect 1875 135 1980 145
rect 2005 215 2045 225
rect 2005 145 2015 215
rect 2035 155 2045 215
rect 2035 145 2085 155
rect 2005 135 2085 145
rect 1895 90 1935 100
rect 1895 70 1905 90
rect 1925 70 1935 90
rect 1895 65 1935 70
rect 1895 45 1905 65
rect 1925 45 1935 65
rect 1895 35 1935 45
rect 1960 75 1980 135
rect 1960 65 2000 75
rect 1960 45 1970 65
rect 1990 45 2000 65
rect 1960 35 2000 45
rect 1810 -65 1820 -45
rect 1840 -65 1850 -45
rect 1750 -130 1790 -120
rect 1450 -160 1490 -150
rect 1750 -150 1760 -130
rect 1780 -150 1790 -130
rect 1750 -160 1790 -150
rect 1390 -260 1400 -190
rect 1420 -260 1430 -190
rect 1390 -270 1430 -260
rect 1470 -190 1510 -180
rect 1470 -260 1480 -190
rect 1500 -260 1510 -190
rect 1470 -270 1510 -260
rect 1535 -190 1575 -180
rect 1535 -260 1545 -190
rect 1565 -260 1575 -190
rect 1535 -270 1575 -260
rect 1600 -190 1640 -180
rect 1600 -260 1610 -190
rect 1630 -260 1640 -190
rect 1600 -270 1640 -260
rect 1665 -190 1705 -180
rect 1665 -260 1675 -190
rect 1695 -260 1705 -190
rect 1665 -270 1705 -260
rect 1730 -190 1770 -180
rect 1730 -260 1740 -190
rect 1760 -260 1770 -190
rect 1730 -270 1770 -260
rect 1810 -190 1850 -65
rect 1875 5 1915 15
rect 1875 -65 1885 5
rect 1905 -65 1915 5
rect 1875 -75 1915 -65
rect 1940 5 1980 15
rect 1940 -65 1950 5
rect 1970 -65 1980 5
rect 1940 -75 1980 -65
rect 2005 5 2045 15
rect 2005 -65 2015 5
rect 2035 -65 2045 5
rect 2005 -75 2045 -65
rect 1960 -105 2000 -95
rect 1960 -125 1970 -105
rect 1990 -125 2000 -105
rect 1960 -135 2000 -125
rect 1960 -180 1980 -135
rect 2065 -180 2085 135
rect 1810 -260 1820 -190
rect 1840 -260 1850 -190
rect 1810 -270 1850 -260
rect 1875 -190 1980 -180
rect 1875 -260 1885 -190
rect 1905 -260 1950 -190
rect 1970 -260 1980 -190
rect 1875 -270 1980 -260
rect 2005 -190 2085 -180
rect 2005 -260 2015 -190
rect 2035 -200 2085 -190
rect 2035 -260 2045 -200
rect 2005 -270 2045 -260
rect 1045 -280 1085 -270
rect 1600 -290 1620 -270
rect 200 -300 240 -290
rect 200 -320 210 -300
rect 230 -310 240 -300
rect 515 -300 620 -290
rect 515 -310 590 -300
rect 230 -320 480 -310
rect 200 -330 480 -320
rect 580 -320 590 -310
rect 610 -320 620 -300
rect 580 -330 620 -320
rect 715 -300 965 -290
rect 1160 -300 1495 -290
rect 715 -320 725 -300
rect 745 -310 1315 -300
rect 745 -320 755 -310
rect 945 -320 1180 -310
rect 1305 -320 1315 -310
rect 1335 -310 1495 -300
rect 1335 -320 1345 -310
rect 715 -330 755 -320
rect 1305 -330 1345 -320
rect 460 -350 480 -330
rect 725 -350 745 -330
rect 460 -370 745 -350
rect 780 -340 820 -330
rect 780 -360 790 -340
rect 810 -350 820 -340
rect 1370 -340 1410 -330
rect 1370 -350 1380 -340
rect 810 -360 1380 -350
rect 1400 -360 1410 -340
rect 780 -370 1410 -360
rect 1475 -350 1495 -310
rect 1515 -300 1620 -290
rect 1515 -320 1525 -300
rect 1545 -310 1620 -300
rect 1830 -300 1870 -290
rect 1545 -320 1555 -310
rect 1515 -330 1555 -320
rect 1830 -320 1840 -300
rect 1860 -320 1870 -300
rect 1830 -330 1870 -320
rect 1830 -350 1850 -330
rect 1475 -370 1850 -350
<< viali >>
rect 210 80 230 90
rect 210 70 230 80
rect 100 -65 120 5
rect 165 -65 185 5
rect 230 -65 250 5
rect 400 145 420 215
rect 610 145 630 215
rect 380 85 400 105
rect 465 65 485 70
rect 465 50 485 65
rect 545 65 565 70
rect 545 50 565 65
rect 680 35 700 55
rect 295 -65 315 -45
rect 100 -260 120 -190
rect 440 -65 460 -45
rect 570 -65 590 -45
rect 885 80 905 100
rect 355 -150 375 -130
rect 715 -65 735 -45
rect 655 -150 675 -130
rect 375 -260 395 -190
rect 440 -260 460 -190
rect 570 -260 590 -190
rect 635 -260 655 -190
rect 780 -65 800 5
rect 845 -65 865 5
rect 1030 145 1050 215
rect 1205 145 1225 215
rect 1505 145 1525 215
rect 1715 145 1735 215
rect 1055 15 1075 85
rect 1105 15 1125 85
rect 1055 -140 1075 -70
rect 1105 -140 1125 -70
rect 1270 -65 1290 5
rect 1335 -65 1355 5
rect 1735 85 1755 105
rect 1435 35 1455 55
rect 1570 65 1590 70
rect 1570 50 1590 65
rect 1650 65 1670 70
rect 1650 50 1670 65
rect 1400 -65 1420 -45
rect 910 -260 930 -190
rect 990 -270 1010 -200
rect 1205 -260 1225 -190
rect 1545 -65 1565 -45
rect 1675 -65 1695 -45
rect 1460 -150 1480 -130
rect 1905 70 1925 90
rect 1820 -65 1840 -45
rect 1760 -150 1780 -130
rect 1480 -260 1500 -190
rect 1545 -260 1565 -190
rect 1675 -260 1695 -190
rect 1740 -260 1760 -190
rect 1885 -65 1905 5
rect 1950 -65 1970 5
rect 2015 -65 2035 5
rect 2015 -260 2035 -190
<< metal1 >>
rect 390 220 430 225
rect 390 140 395 220
rect 425 140 430 220
rect 390 135 430 140
rect 600 220 640 225
rect 600 140 605 220
rect 635 140 640 220
rect 1020 215 1060 225
rect 1020 150 1030 215
rect 600 135 640 140
rect 900 145 1030 150
rect 1050 145 1060 215
rect 900 135 1060 145
rect 1195 215 1235 225
rect 1195 145 1205 215
rect 1225 145 1235 215
rect 1195 135 1235 145
rect 1495 220 1535 225
rect 1495 140 1500 220
rect 1530 140 1535 220
rect 1495 135 1535 140
rect 1705 220 1745 225
rect 1705 140 1710 220
rect 1740 140 1745 220
rect 1705 135 1745 140
rect 370 105 410 115
rect 900 110 915 135
rect 200 90 240 100
rect 200 70 210 90
rect 230 70 240 90
rect 370 85 380 105
rect 400 85 410 105
rect 875 100 915 110
rect 370 75 410 85
rect 640 80 850 95
rect 200 60 240 70
rect 115 30 290 45
rect 115 15 130 30
rect 90 5 130 15
rect 90 -65 100 5
rect 120 -65 130 5
rect 90 -75 130 -65
rect 155 5 195 15
rect 155 -65 165 5
rect 185 -65 195 5
rect 155 -75 195 -65
rect 220 10 260 15
rect 220 -70 225 10
rect 255 -70 260 10
rect 275 -5 290 30
rect 395 25 410 75
rect 455 70 495 80
rect 455 50 465 70
rect 485 50 495 70
rect 455 40 495 50
rect 535 70 575 80
rect 535 50 545 70
rect 565 50 575 70
rect 535 40 575 50
rect 640 25 655 80
rect 670 55 710 65
rect 670 35 680 55
rect 700 35 710 55
rect 670 25 710 35
rect 395 10 655 25
rect 675 -5 690 25
rect 835 15 850 80
rect 875 80 885 100
rect 905 80 915 100
rect 875 70 915 80
rect 275 -20 690 -5
rect 770 5 810 15
rect 220 -75 260 -70
rect 285 -45 470 -35
rect 285 -65 295 -45
rect 315 -65 440 -45
rect 460 -65 470 -45
rect 285 -75 470 -65
rect 560 -45 745 -35
rect 560 -65 570 -45
rect 590 -65 715 -45
rect 735 -65 745 -45
rect 560 -75 745 -65
rect 770 -65 780 5
rect 800 -65 810 5
rect 770 -75 810 -65
rect 835 5 875 15
rect 835 -65 845 5
rect 865 -65 875 5
rect 835 -75 875 -65
rect 180 -90 195 -75
rect 770 -90 785 -75
rect 180 -105 785 -90
rect 345 -130 385 -120
rect 345 -150 355 -130
rect 375 -140 385 -130
rect 645 -130 685 -120
rect 645 -140 655 -130
rect 375 -150 450 -140
rect 345 -160 450 -150
rect 430 -180 450 -160
rect 580 -150 655 -140
rect 675 -150 685 -130
rect 580 -160 685 -150
rect 580 -180 600 -160
rect 90 -190 130 -180
rect 90 -260 100 -190
rect 120 -260 130 -190
rect 90 -270 130 -260
rect 365 -185 405 -180
rect 365 -265 370 -185
rect 400 -265 405 -185
rect 365 -270 405 -265
rect 430 -190 470 -180
rect 430 -260 440 -190
rect 460 -260 470 -190
rect 430 -270 470 -260
rect 560 -190 600 -180
rect 560 -260 570 -190
rect 590 -260 600 -190
rect 560 -270 600 -260
rect 625 -185 665 -180
rect 625 -265 630 -185
rect 660 -265 665 -185
rect 625 -270 665 -265
rect 900 -190 940 -180
rect 900 -260 910 -190
rect 930 -260 940 -190
rect 900 -270 940 -260
rect 980 -190 995 135
rect 1045 90 1135 95
rect 1045 10 1050 90
rect 1080 10 1100 90
rect 1130 10 1135 90
rect 1045 5 1135 10
rect 1045 -65 1135 -60
rect 1045 -145 1050 -65
rect 1080 -145 1100 -65
rect 1130 -145 1135 -65
rect 1045 -150 1135 -145
rect 1220 -180 1235 135
rect 1725 105 1765 115
rect 1285 80 1495 95
rect 1725 85 1735 105
rect 1755 85 1765 105
rect 1285 15 1300 80
rect 1425 55 1465 65
rect 1425 35 1435 55
rect 1455 35 1465 55
rect 1425 25 1465 35
rect 1480 25 1495 80
rect 1560 70 1600 80
rect 1560 50 1570 70
rect 1590 50 1600 70
rect 1560 40 1600 50
rect 1640 70 1680 80
rect 1640 50 1650 70
rect 1670 50 1680 70
rect 1640 40 1680 50
rect 1725 75 1765 85
rect 1895 90 1935 100
rect 1725 25 1740 75
rect 1895 70 1905 90
rect 1925 70 1935 90
rect 1895 60 1935 70
rect 1260 5 1300 15
rect 1260 -65 1270 5
rect 1290 -65 1300 5
rect 1260 -75 1300 -65
rect 1325 5 1365 15
rect 1325 -65 1335 5
rect 1355 -65 1365 5
rect 1445 -5 1460 25
rect 1480 10 1740 25
rect 1845 30 2020 45
rect 1845 -5 1860 30
rect 2005 15 2020 30
rect 1445 -20 1860 -5
rect 1875 10 1915 15
rect 1325 -75 1365 -65
rect 1390 -45 1575 -35
rect 1390 -65 1400 -45
rect 1420 -65 1545 -45
rect 1565 -65 1575 -45
rect 1390 -75 1575 -65
rect 1665 -45 1850 -35
rect 1665 -65 1675 -45
rect 1695 -65 1820 -45
rect 1840 -65 1850 -45
rect 1665 -75 1850 -65
rect 1875 -70 1880 10
rect 1910 -70 1915 10
rect 1875 -75 1915 -70
rect 1940 5 1980 15
rect 1940 -65 1950 5
rect 1970 -65 1980 5
rect 1940 -75 1980 -65
rect 2005 5 2045 15
rect 2005 -65 2015 5
rect 2035 -65 2045 5
rect 2005 -75 2045 -65
rect 1350 -90 1365 -75
rect 1940 -90 1955 -75
rect 1350 -105 1955 -90
rect 1450 -130 1490 -120
rect 1450 -150 1460 -130
rect 1480 -140 1490 -130
rect 1750 -130 1790 -120
rect 1750 -140 1760 -130
rect 1480 -150 1555 -140
rect 1450 -160 1555 -150
rect 1535 -180 1555 -160
rect 1685 -150 1760 -140
rect 1780 -150 1790 -130
rect 1685 -160 1790 -150
rect 1685 -180 1705 -160
rect 1195 -190 1235 -180
rect 980 -200 1020 -190
rect 980 -270 990 -200
rect 1010 -270 1020 -200
rect 1195 -260 1205 -190
rect 1225 -260 1235 -190
rect 1195 -270 1235 -260
rect 1470 -185 1510 -180
rect 1470 -265 1475 -185
rect 1505 -265 1510 -185
rect 1470 -270 1510 -265
rect 1535 -190 1575 -180
rect 1535 -260 1545 -190
rect 1565 -260 1575 -190
rect 1535 -270 1575 -260
rect 1665 -190 1705 -180
rect 1665 -260 1675 -190
rect 1695 -260 1705 -190
rect 1665 -270 1705 -260
rect 1730 -185 1770 -180
rect 1730 -265 1735 -185
rect 1765 -265 1770 -185
rect 1730 -270 1770 -265
rect 2005 -190 2045 -180
rect 2005 -260 2015 -190
rect 2035 -260 2045 -190
rect 2005 -270 2045 -260
rect 115 -285 130 -270
rect 900 -285 915 -270
rect 980 -280 1020 -270
rect 115 -300 915 -285
rect 1220 -285 1235 -270
rect 2005 -285 2020 -270
rect 1220 -300 2020 -285
<< via1 >>
rect 395 215 425 220
rect 395 145 400 215
rect 400 145 420 215
rect 420 145 425 215
rect 395 140 425 145
rect 605 215 635 220
rect 605 145 610 215
rect 610 145 630 215
rect 630 145 635 215
rect 605 140 635 145
rect 1500 215 1530 220
rect 1500 145 1505 215
rect 1505 145 1525 215
rect 1525 145 1530 215
rect 1500 140 1530 145
rect 1710 215 1740 220
rect 1710 145 1715 215
rect 1715 145 1735 215
rect 1735 145 1740 215
rect 1710 140 1740 145
rect 225 5 255 10
rect 225 -65 230 5
rect 230 -65 250 5
rect 250 -65 255 5
rect 225 -70 255 -65
rect 370 -190 400 -185
rect 370 -260 375 -190
rect 375 -260 395 -190
rect 395 -260 400 -190
rect 370 -265 400 -260
rect 630 -190 660 -185
rect 630 -260 635 -190
rect 635 -260 655 -190
rect 655 -260 660 -190
rect 630 -265 660 -260
rect 1050 85 1080 90
rect 1050 15 1055 85
rect 1055 15 1075 85
rect 1075 15 1080 85
rect 1050 10 1080 15
rect 1100 85 1130 90
rect 1100 15 1105 85
rect 1105 15 1125 85
rect 1125 15 1130 85
rect 1100 10 1130 15
rect 1050 -70 1080 -65
rect 1050 -140 1055 -70
rect 1055 -140 1075 -70
rect 1075 -140 1080 -70
rect 1050 -145 1080 -140
rect 1100 -70 1130 -65
rect 1100 -140 1105 -70
rect 1105 -140 1125 -70
rect 1125 -140 1130 -70
rect 1100 -145 1130 -140
rect 1880 5 1910 10
rect 1880 -65 1885 5
rect 1885 -65 1905 5
rect 1905 -65 1910 5
rect 1880 -70 1910 -65
rect 1475 -190 1505 -185
rect 1475 -260 1480 -190
rect 1480 -260 1500 -190
rect 1500 -260 1505 -190
rect 1475 -265 1505 -260
rect 1735 -190 1765 -185
rect 1735 -260 1740 -190
rect 1740 -260 1760 -190
rect 1760 -260 1765 -190
rect 1735 -265 1765 -260
<< metal2 >>
rect 390 220 1745 225
rect 390 140 395 220
rect 425 140 605 220
rect 635 140 1500 220
rect 1530 140 1710 220
rect 1740 140 1745 220
rect 390 135 1745 140
rect 1045 90 1135 135
rect 220 10 260 15
rect 220 -70 225 10
rect 255 -70 260 10
rect 1045 10 1050 90
rect 1080 10 1100 90
rect 1130 10 1135 90
rect 1045 5 1135 10
rect 1875 10 1915 15
rect 220 -180 260 -70
rect 1045 -65 1135 -60
rect 1045 -145 1050 -65
rect 1080 -145 1100 -65
rect 1130 -145 1135 -65
rect 1045 -180 1135 -145
rect 1875 -70 1880 10
rect 1910 -70 1915 10
rect 1875 -180 1915 -70
rect 220 -185 1915 -180
rect 220 -265 370 -185
rect 400 -265 630 -185
rect 660 -265 1475 -185
rect 1505 -265 1735 -185
rect 1765 -265 1915 -185
rect 220 -270 1915 -265
<< labels >>
rlabel poly 1030 -300 1030 -300 5 SH
rlabel poly 1070 260 1070 260 1 Shb
rlabel locali 915 90 915 90 3 C-
rlabel locali 1220 70 1220 70 7 C+
<< end >>
