magic
tech sky130A
timestamp 1702648776
<< nwell >>
rect 170 2170 345 2310
<< nmos >>
rect 240 2035 255 2135
<< pmos >>
rect 240 2190 255 2290
<< ndiff >>
rect 190 2120 240 2135
rect 190 2050 205 2120
rect 225 2050 240 2120
rect 190 2035 240 2050
rect 255 2120 305 2135
rect 255 2050 270 2120
rect 290 2050 305 2120
rect 255 2035 305 2050
<< pdiff >>
rect 190 2275 240 2290
rect 190 2205 205 2275
rect 225 2205 240 2275
rect 190 2190 240 2205
rect 255 2275 305 2290
rect 255 2205 270 2275
rect 290 2205 305 2275
rect 255 2190 305 2205
<< ndiffc >>
rect 205 2050 225 2120
rect 270 2050 290 2120
<< pdiffc >>
rect 205 2205 225 2275
rect 270 2205 290 2275
<< poly >>
rect 280 2335 320 2345
rect 280 2315 290 2335
rect 310 2320 320 2335
rect 310 2315 405 2320
rect 280 2305 405 2315
rect 240 2290 255 2305
rect 240 2135 255 2190
rect 240 1665 255 2035
rect 240 1650 420 1665
<< polycont >>
rect 290 2315 310 2335
<< locali >>
rect 280 2335 320 2345
rect 280 2315 290 2335
rect 310 2315 320 2335
rect 280 2305 320 2315
rect 280 2285 300 2305
rect 195 2275 235 2285
rect 195 2205 205 2275
rect 225 2205 235 2275
rect 195 2195 235 2205
rect 260 2275 300 2285
rect 260 2205 270 2275
rect 290 2205 300 2275
rect 195 2120 235 2130
rect 195 2050 205 2120
rect 225 2050 235 2120
rect 195 2040 235 2050
rect 260 2120 300 2205
rect 260 2050 270 2120
rect 290 2050 300 2120
rect 260 2040 300 2050
rect 2350 810 2390 820
rect 2350 790 2360 810
rect 2380 790 2390 810
rect 2350 780 2390 790
<< viali >>
rect 1690 2315 1710 2335
rect 205 2205 225 2275
rect 205 2050 225 2120
rect 300 1595 320 1615
rect 2360 1600 2380 1620
rect 2360 790 2380 810
<< metal1 >>
rect 1680 2340 1720 2345
rect 1680 2310 1685 2340
rect 1715 2310 1720 2340
rect 1680 2305 1720 2310
rect 2230 2340 2445 2345
rect 2230 2310 2235 2340
rect 2265 2310 2445 2340
rect 2230 2305 2445 2310
rect 195 2280 235 2285
rect 195 2200 200 2280
rect 230 2200 235 2280
rect 195 2195 235 2200
rect 195 2125 235 2130
rect 195 2045 200 2125
rect 230 2045 235 2125
rect 195 2040 235 2045
rect 290 2120 510 2160
rect 2165 2120 2390 2160
rect 290 1615 330 2120
rect 290 1595 300 1615
rect 320 1595 330 1615
rect 290 1585 330 1595
rect 2350 1620 2390 2120
rect 2405 1680 2445 2305
rect 2405 1640 2645 1680
rect 2350 1600 2360 1620
rect 2380 1600 2390 1620
rect 2350 1590 2390 1600
rect 2605 820 2645 1640
rect 2350 810 2645 820
rect 2350 790 2360 810
rect 2380 790 2645 810
rect 2350 780 2645 790
<< via1 >>
rect 1685 2335 1715 2340
rect 1685 2315 1690 2335
rect 1690 2315 1710 2335
rect 1710 2315 1715 2335
rect 1685 2310 1715 2315
rect 2235 2310 2265 2340
rect 200 2275 230 2280
rect 200 2205 205 2275
rect 205 2205 225 2275
rect 225 2205 230 2275
rect 200 2200 230 2205
rect 200 2120 230 2125
rect 200 2050 205 2120
rect 205 2050 225 2120
rect 225 2050 230 2120
rect 200 2045 230 2050
<< metal2 >>
rect 1680 2340 2270 2345
rect 1680 2310 1685 2340
rect 1715 2310 2235 2340
rect 2265 2310 2270 2340
rect 1680 2305 2270 2310
rect 195 2280 665 2285
rect 195 2200 200 2280
rect 230 2200 665 2280
rect 195 2195 665 2200
rect 2015 2195 2390 2285
rect 195 2125 530 2135
rect 195 2045 200 2125
rect 230 2045 530 2125
rect 195 1880 530 2045
rect 0 1790 560 1880
rect 0 0 45 1790
rect 2350 1630 2390 2195
use bias_cg  bias_cg_0
timestamp 1702648396
transform 1 0 385 0 1 970
box -385 -970 2311 660
use middle  middle_0
timestamp 1702643716
transform 1 0 270 0 1 2060
box 50 -410 2085 405
<< end >>
