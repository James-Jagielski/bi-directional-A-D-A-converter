magic
tech sky130A
magscale 1 2
timestamp 1702589910
<< nwell >>
rect -180 660 1240 1430
<< nmos >>
rect -40 300 -10 500
rect 90 300 120 500
rect 220 300 250 500
rect 350 300 380 500
rect 480 300 510 500
rect 770 300 800 500
rect -40 -330 -10 -130
rect 90 -330 120 -130
rect 220 -330 250 -130
rect 350 -330 380 -130
rect 480 -330 510 -130
rect 610 -330 640 -130
rect 740 -330 770 -130
<< pmos >>
rect -40 770 -10 970
rect 40 770 70 970
rect 170 770 200 970
rect 460 770 490 970
rect 590 770 620 970
rect 670 770 700 970
rect 960 770 990 970
<< ndiff >>
rect -140 470 -40 500
rect -140 330 -110 470
rect -70 330 -40 470
rect -140 300 -40 330
rect -10 470 90 500
rect -10 330 20 470
rect 60 330 90 470
rect -10 300 90 330
rect 120 470 220 500
rect 120 330 150 470
rect 190 330 220 470
rect 120 300 220 330
rect 250 470 350 500
rect 250 330 280 470
rect 320 330 350 470
rect 250 300 350 330
rect 380 470 480 500
rect 380 330 410 470
rect 450 330 480 470
rect 380 300 480 330
rect 510 470 610 500
rect 510 330 540 470
rect 580 330 610 470
rect 510 300 610 330
rect 670 470 770 500
rect 670 330 700 470
rect 740 330 770 470
rect 670 300 770 330
rect 800 470 900 500
rect 800 330 830 470
rect 870 330 900 470
rect 800 300 900 330
rect -140 -160 -40 -130
rect -140 -300 -110 -160
rect -70 -300 -40 -160
rect -140 -330 -40 -300
rect -10 -160 90 -130
rect -10 -300 20 -160
rect 60 -300 90 -160
rect -10 -330 90 -300
rect 120 -160 220 -130
rect 120 -300 150 -160
rect 190 -300 220 -160
rect 120 -330 220 -300
rect 250 -160 350 -130
rect 250 -300 280 -160
rect 320 -300 350 -160
rect 250 -330 350 -300
rect 380 -160 480 -130
rect 380 -300 410 -160
rect 450 -300 480 -160
rect 380 -330 480 -300
rect 510 -160 610 -130
rect 510 -300 540 -160
rect 580 -300 610 -160
rect 510 -330 610 -300
rect 640 -160 740 -130
rect 640 -300 670 -160
rect 710 -300 740 -160
rect 640 -330 740 -300
rect 770 -160 870 -130
rect 770 -300 800 -160
rect 840 -300 870 -160
rect 770 -330 870 -300
<< pdiff >>
rect -140 940 -40 970
rect -140 800 -110 940
rect -70 800 -40 940
rect -140 770 -40 800
rect -10 770 40 970
rect 70 940 170 970
rect 70 800 100 940
rect 140 800 170 940
rect 70 770 170 800
rect 200 940 300 970
rect 200 800 230 940
rect 270 800 300 940
rect 200 770 300 800
rect 360 940 460 970
rect 360 800 390 940
rect 430 800 460 940
rect 360 770 460 800
rect 490 940 590 970
rect 490 800 520 940
rect 560 800 590 940
rect 490 770 590 800
rect 620 770 670 970
rect 700 940 800 970
rect 700 800 730 940
rect 770 800 800 940
rect 700 770 800 800
rect 860 940 960 970
rect 860 800 890 940
rect 930 800 960 940
rect 860 770 960 800
rect 990 940 1090 970
rect 990 800 1020 940
rect 1060 800 1090 940
rect 990 770 1090 800
<< ndiffc >>
rect -110 330 -70 470
rect 20 330 60 470
rect 150 330 190 470
rect 280 330 320 470
rect 410 330 450 470
rect 540 330 580 470
rect 700 330 740 470
rect 830 330 870 470
rect -110 -300 -70 -160
rect 20 -300 60 -160
rect 150 -300 190 -160
rect 280 -300 320 -160
rect 410 -300 450 -160
rect 540 -300 580 -160
rect 670 -300 710 -160
rect 800 -300 840 -160
<< pdiffc >>
rect -110 800 -70 940
rect 100 800 140 940
rect 230 800 270 940
rect 390 800 430 940
rect 520 800 560 940
rect 730 800 770 940
rect 890 800 930 940
rect 1020 800 1060 940
<< psubdiff >>
rect -210 -620 1250 -590
rect -210 -760 -180 -620
rect -140 -760 -100 -620
rect -60 -760 -20 -620
rect 20 -760 60 -620
rect 100 -760 140 -620
rect 180 -760 220 -620
rect 260 -760 300 -620
rect 340 -760 380 -620
rect 420 -760 460 -620
rect 500 -760 540 -620
rect 580 -760 620 -620
rect 660 -760 700 -620
rect 740 -760 780 -620
rect 820 -760 860 -620
rect 900 -760 940 -620
rect 980 -760 1020 -620
rect 1060 -760 1100 -620
rect 1140 -760 1180 -620
rect 1220 -760 1250 -620
rect -210 -790 1250 -760
<< nsubdiff >>
rect -140 1360 1110 1390
rect -140 1220 -110 1360
rect -70 1220 -30 1360
rect 10 1220 50 1360
rect 90 1220 130 1360
rect 170 1220 210 1360
rect 250 1220 290 1360
rect 330 1220 370 1360
rect 410 1220 450 1360
rect 490 1220 530 1360
rect 570 1220 610 1360
rect 650 1220 690 1360
rect 730 1220 770 1360
rect 810 1220 850 1360
rect 890 1220 930 1360
rect 970 1220 1010 1360
rect 1050 1220 1110 1360
rect -140 1190 1110 1220
<< psubdiffcont >>
rect -180 -760 -140 -620
rect -100 -760 -60 -620
rect -20 -760 20 -620
rect 60 -760 100 -620
rect 140 -760 180 -620
rect 220 -760 260 -620
rect 300 -760 340 -620
rect 380 -760 420 -620
rect 460 -760 500 -620
rect 540 -760 580 -620
rect 620 -760 660 -620
rect 700 -760 740 -620
rect 780 -760 820 -620
rect 860 -760 900 -620
rect 940 -760 980 -620
rect 1020 -760 1060 -620
rect 1100 -760 1140 -620
rect 1180 -760 1220 -620
<< nsubdiffcont >>
rect -110 1220 -70 1360
rect -30 1220 10 1360
rect 50 1220 90 1360
rect 130 1220 170 1360
rect 210 1220 250 1360
rect 290 1220 330 1360
rect 370 1220 410 1360
rect 450 1220 490 1360
rect 530 1220 570 1360
rect 610 1220 650 1360
rect 690 1220 730 1360
rect 770 1220 810 1360
rect 850 1220 890 1360
rect 930 1220 970 1360
rect 1010 1220 1050 1360
<< poly >>
rect 200 1060 280 1080
rect 200 1030 220 1060
rect 40 1020 220 1030
rect 260 1020 280 1060
rect 40 1000 280 1020
rect 380 1060 460 1080
rect 380 1020 400 1060
rect 440 1030 460 1060
rect 670 1050 1280 1080
rect 440 1020 620 1030
rect 380 1000 620 1020
rect -40 970 -10 1000
rect 40 970 70 1000
rect 170 970 200 1000
rect 460 970 490 1000
rect 590 970 620 1000
rect 670 970 700 1050
rect 960 970 990 1000
rect -40 690 -10 770
rect 40 740 70 770
rect 170 740 200 770
rect 460 740 490 770
rect 590 740 620 770
rect 670 690 700 770
rect -270 660 700 690
rect 960 740 990 770
rect 960 710 1280 740
rect 90 580 510 610
rect 90 560 120 580
rect -270 530 120 560
rect -40 500 -10 530
rect 90 500 120 530
rect 220 500 250 530
rect 350 500 380 530
rect 480 500 510 580
rect 770 500 800 530
rect -40 270 -10 300
rect 90 270 120 300
rect 220 220 250 300
rect -270 190 250 220
rect 350 140 380 300
rect 480 270 510 300
rect 770 270 800 300
rect 960 270 990 710
rect 770 250 850 270
rect 770 210 790 250
rect 830 210 850 250
rect 770 190 850 210
rect 910 250 990 270
rect 910 210 930 250
rect 970 210 990 250
rect 910 190 990 210
rect 350 110 1290 140
rect 90 40 970 60
rect 90 30 910 40
rect -270 -100 -10 -70
rect -40 -130 -10 -100
rect 90 -130 120 30
rect 350 -40 430 -20
rect 350 -80 370 -40
rect 410 -80 430 -40
rect 350 -100 430 -80
rect 600 -40 680 -20
rect 600 -80 620 -40
rect 660 -80 680 -40
rect 600 -100 680 -80
rect 220 -130 250 -100
rect 350 -130 380 -100
rect 480 -130 510 -100
rect 610 -130 640 -100
rect 740 -130 770 30
rect 890 0 910 30
rect 950 0 970 40
rect 890 -20 970 0
rect -40 -360 -10 -330
rect 90 -360 120 -330
rect 220 -490 250 -330
rect 350 -360 380 -330
rect 300 -380 380 -360
rect 300 -420 320 -380
rect 360 -420 380 -380
rect 300 -440 380 -420
rect 480 -360 510 -330
rect 610 -360 640 -330
rect 740 -360 770 -330
rect 480 -380 560 -360
rect 480 -420 500 -380
rect 540 -420 560 -380
rect 480 -440 560 -420
rect 220 -520 1290 -490
<< polycont >>
rect 220 1020 260 1060
rect 400 1020 440 1060
rect 790 210 830 250
rect 930 210 970 250
rect 370 -80 410 -40
rect 620 -80 660 -40
rect 910 0 950 40
rect 320 -420 360 -380
rect 500 -420 540 -380
<< locali >>
rect -130 1360 1100 1380
rect -130 1220 -110 1360
rect -70 1220 -30 1360
rect 10 1220 50 1360
rect 90 1220 130 1360
rect 170 1220 210 1360
rect 250 1220 290 1360
rect 330 1220 370 1360
rect 410 1220 450 1360
rect 490 1220 530 1360
rect 570 1220 610 1360
rect 650 1220 690 1360
rect 730 1220 770 1360
rect 810 1220 850 1360
rect 890 1220 930 1360
rect 970 1220 1010 1360
rect 1050 1220 1100 1360
rect -130 1200 1100 1220
rect 1150 1180 1230 1200
rect 1150 1160 1170 1180
rect -90 1140 1170 1160
rect 1210 1160 1230 1180
rect 1210 1140 1280 1160
rect -90 1120 1280 1140
rect -90 960 -50 1120
rect 200 1060 280 1080
rect 200 1020 220 1060
rect 260 1020 280 1060
rect 200 1000 280 1020
rect 380 1060 460 1080
rect 380 1020 400 1060
rect 440 1020 460 1060
rect 380 1000 460 1020
rect 750 1000 1280 1040
rect 210 960 250 1000
rect 410 960 450 1000
rect 750 960 790 1000
rect -130 940 -50 960
rect -130 800 -110 940
rect -70 800 -50 940
rect -130 780 -50 800
rect 80 940 160 960
rect 80 800 100 940
rect 140 800 160 940
rect 80 780 160 800
rect 210 940 290 960
rect 210 800 230 940
rect 270 800 290 940
rect 210 780 290 800
rect 250 720 290 780
rect 170 680 290 720
rect 370 940 450 960
rect 370 800 390 940
rect 430 800 450 940
rect 370 780 450 800
rect 500 940 580 960
rect 500 800 520 940
rect 560 800 580 940
rect 500 780 580 800
rect 710 940 790 960
rect 710 800 730 940
rect 770 800 790 940
rect 710 780 790 800
rect 870 940 950 960
rect 870 800 890 940
rect 930 800 950 940
rect 870 780 950 800
rect 1000 940 1080 960
rect 1000 800 1020 940
rect 1060 800 1080 940
rect 1000 780 1080 800
rect 370 720 410 780
rect 750 750 790 780
rect 370 680 430 720
rect 750 710 850 750
rect 170 490 210 680
rect 390 490 430 680
rect 810 490 850 710
rect -130 470 -50 490
rect -130 330 -110 470
rect -70 330 -50 470
rect -130 310 -50 330
rect 0 470 80 490
rect 0 330 20 470
rect 60 330 80 470
rect 0 310 80 330
rect 130 470 210 490
rect 130 330 150 470
rect 190 330 210 470
rect 130 310 210 330
rect 260 470 340 490
rect 260 330 280 470
rect 320 330 340 470
rect 260 310 340 330
rect 390 470 470 490
rect 390 330 410 470
rect 450 330 470 470
rect 390 310 470 330
rect 520 470 600 490
rect 520 330 540 470
rect 580 330 600 470
rect 520 310 600 330
rect 680 470 760 490
rect 680 330 700 470
rect 740 330 760 470
rect 680 310 760 330
rect 810 470 890 490
rect 810 330 830 470
rect 870 330 890 470
rect 810 310 890 330
rect -90 270 -50 310
rect 260 270 300 310
rect -90 230 300 270
rect 680 80 720 310
rect 770 250 850 270
rect 770 210 790 250
rect 830 210 850 250
rect 770 190 850 210
rect 910 250 990 270
rect 910 210 930 250
rect 970 210 990 250
rect 910 190 990 210
rect 260 40 720 80
rect 260 -140 300 40
rect 350 -40 430 -20
rect 350 -80 370 -40
rect 410 -60 430 -40
rect 600 -40 680 -20
rect 410 -80 560 -60
rect 350 -100 560 -80
rect 600 -80 620 -40
rect 660 -60 680 -40
rect 780 -60 820 190
rect 930 60 970 190
rect 890 40 970 60
rect 890 0 910 40
rect 950 0 970 40
rect 890 -20 970 0
rect 1040 -60 1080 780
rect 660 -80 1080 -60
rect 600 -100 1080 -80
rect 1160 930 1240 950
rect 1160 890 1180 930
rect 1220 890 1240 930
rect 1160 870 1240 890
rect 520 -140 560 -100
rect 780 -140 820 -100
rect -130 -160 -50 -140
rect -130 -300 -110 -160
rect -70 -300 -50 -160
rect -130 -340 -50 -300
rect 0 -160 80 -140
rect 0 -300 20 -160
rect 60 -300 80 -160
rect 0 -320 80 -300
rect -130 -380 -110 -340
rect -70 -380 -50 -340
rect -130 -400 -50 -380
rect -90 -520 -50 -400
rect 40 -440 80 -320
rect 130 -160 210 -140
rect 130 -300 150 -160
rect 190 -300 210 -160
rect 130 -340 210 -300
rect 260 -160 340 -140
rect 260 -300 280 -160
rect 320 -300 340 -160
rect 260 -320 340 -300
rect 390 -160 470 -140
rect 390 -300 410 -160
rect 450 -300 470 -160
rect 390 -320 470 -300
rect 520 -160 600 -140
rect 520 -300 540 -160
rect 580 -300 600 -160
rect 520 -320 600 -300
rect 650 -160 730 -140
rect 650 -300 670 -160
rect 710 -300 730 -160
rect 650 -320 730 -300
rect 780 -160 860 -140
rect 780 -300 800 -160
rect 840 -300 860 -160
rect 780 -320 860 -300
rect 130 -380 150 -340
rect 190 -380 210 -340
rect 690 -360 730 -320
rect 1160 -360 1200 870
rect 130 -400 210 -380
rect 300 -380 380 -360
rect 300 -420 320 -380
rect 360 -420 380 -380
rect 300 -440 380 -420
rect 480 -380 560 -360
rect 480 -420 500 -380
rect 540 -420 560 -380
rect 690 -400 1200 -360
rect 480 -440 560 -420
rect 40 -480 340 -440
rect 480 -520 520 -440
rect -90 -560 520 -520
rect -200 -620 1240 -600
rect -200 -760 -180 -620
rect -140 -760 -100 -620
rect -60 -760 -20 -620
rect 20 -760 60 -620
rect 100 -760 140 -620
rect 180 -760 220 -620
rect 260 -760 300 -620
rect 340 -760 380 -620
rect 420 -760 460 -620
rect 500 -760 540 -620
rect 580 -760 620 -620
rect 660 -760 700 -620
rect 740 -760 780 -620
rect 820 -760 860 -620
rect 900 -760 940 -620
rect 980 -760 1020 -620
rect 1060 -760 1100 -620
rect 1140 -760 1180 -620
rect 1220 -760 1240 -620
rect -200 -780 1240 -760
<< viali >>
rect -110 1220 -70 1360
rect -30 1220 10 1360
rect 50 1220 90 1360
rect 130 1220 170 1360
rect 210 1220 250 1360
rect 290 1220 330 1360
rect 370 1220 410 1360
rect 450 1220 490 1360
rect 530 1220 570 1360
rect 610 1220 650 1360
rect 690 1220 730 1360
rect 770 1220 810 1360
rect 850 1220 890 1360
rect 930 1220 970 1360
rect 1010 1220 1050 1360
rect 1170 1140 1210 1180
rect 100 800 140 940
rect 520 800 560 940
rect 890 800 930 940
rect 20 330 60 470
rect 540 330 580 470
rect 1180 890 1220 930
rect -110 -380 -70 -340
rect 410 -300 450 -160
rect 150 -380 190 -340
rect -180 -760 -140 -620
rect -100 -760 -60 -620
rect -20 -760 20 -620
rect 60 -760 100 -620
rect 140 -760 180 -620
rect 220 -760 260 -620
rect 300 -760 340 -620
rect 380 -760 420 -620
rect 460 -760 500 -620
rect 540 -760 580 -620
rect 620 -760 660 -620
rect 700 -760 740 -620
rect 780 -760 820 -620
rect 860 -760 900 -620
rect 940 -760 980 -620
rect 1020 -760 1060 -620
rect 1100 -760 1140 -620
rect 1180 -760 1220 -620
<< metal1 >>
rect -130 1370 1100 1380
rect -130 1210 -120 1370
rect 1090 1210 1100 1370
rect -130 1200 1100 1210
rect 1150 1180 1230 1200
rect 1150 1140 1170 1180
rect 1210 1140 1230 1180
rect 1150 1120 1230 1140
rect 80 950 160 960
rect 80 790 90 950
rect 150 790 160 950
rect 80 780 160 790
rect 500 950 580 960
rect 500 790 510 950
rect 570 790 580 950
rect 500 780 580 790
rect 870 950 950 960
rect 870 790 880 950
rect 940 790 950 950
rect 1160 950 1200 1120
rect 1160 930 1240 950
rect 1160 890 1180 930
rect 1220 890 1240 930
rect 1160 870 1240 890
rect 870 780 950 790
rect 0 480 80 500
rect 0 320 10 480
rect 70 320 80 480
rect 0 300 80 320
rect 510 480 610 500
rect 510 320 530 480
rect 590 320 610 480
rect 510 300 610 320
rect 380 -150 480 -130
rect 380 -310 400 -150
rect 460 -310 480 -150
rect -130 -340 210 -320
rect 380 -330 480 -310
rect -130 -380 -110 -340
rect -70 -380 150 -340
rect 190 -380 210 -340
rect -130 -400 210 -380
rect -210 -610 1250 -590
rect -210 -770 -190 -610
rect 1230 -770 1250 -610
rect -210 -790 1250 -770
<< via1 >>
rect -120 1360 1090 1370
rect -120 1220 -110 1360
rect -110 1220 -70 1360
rect -70 1220 -30 1360
rect -30 1220 10 1360
rect 10 1220 50 1360
rect 50 1220 90 1360
rect 90 1220 130 1360
rect 130 1220 170 1360
rect 170 1220 210 1360
rect 210 1220 250 1360
rect 250 1220 290 1360
rect 290 1220 330 1360
rect 330 1220 370 1360
rect 370 1220 410 1360
rect 410 1220 450 1360
rect 450 1220 490 1360
rect 490 1220 530 1360
rect 530 1220 570 1360
rect 570 1220 610 1360
rect 610 1220 650 1360
rect 650 1220 690 1360
rect 690 1220 730 1360
rect 730 1220 770 1360
rect 770 1220 810 1360
rect 810 1220 850 1360
rect 850 1220 890 1360
rect 890 1220 930 1360
rect 930 1220 970 1360
rect 970 1220 1010 1360
rect 1010 1220 1050 1360
rect 1050 1220 1090 1360
rect -120 1210 1090 1220
rect 90 940 150 950
rect 90 800 100 940
rect 100 800 140 940
rect 140 800 150 940
rect 90 790 150 800
rect 510 940 570 950
rect 510 800 520 940
rect 520 800 560 940
rect 560 800 570 940
rect 510 790 570 800
rect 880 940 940 950
rect 880 800 890 940
rect 890 800 930 940
rect 930 800 940 940
rect 880 790 940 800
rect 10 470 70 480
rect 10 330 20 470
rect 20 330 60 470
rect 60 330 70 470
rect 10 320 70 330
rect 530 470 590 480
rect 530 330 540 470
rect 540 330 580 470
rect 580 330 590 470
rect 530 320 590 330
rect 400 -160 460 -150
rect 400 -300 410 -160
rect 410 -300 450 -160
rect 450 -300 460 -160
rect 400 -310 460 -300
rect -190 -620 1230 -610
rect -190 -760 -180 -620
rect -180 -760 -140 -620
rect -140 -760 -100 -620
rect -100 -760 -60 -620
rect -60 -760 -20 -620
rect -20 -760 20 -620
rect 20 -760 60 -620
rect 60 -760 100 -620
rect 100 -760 140 -620
rect 140 -760 180 -620
rect 180 -760 220 -620
rect 220 -760 260 -620
rect 260 -760 300 -620
rect 300 -760 340 -620
rect 340 -760 380 -620
rect 380 -760 420 -620
rect 420 -760 460 -620
rect 460 -760 500 -620
rect 500 -760 540 -620
rect 540 -760 580 -620
rect 580 -760 620 -620
rect 620 -760 660 -620
rect 660 -760 700 -620
rect 700 -760 740 -620
rect 740 -760 780 -620
rect 780 -760 820 -620
rect 820 -760 860 -620
rect 860 -760 900 -620
rect 900 -760 940 -620
rect 940 -760 980 -620
rect 980 -760 1020 -620
rect 1020 -760 1060 -620
rect 1060 -760 1100 -620
rect 1100 -760 1140 -620
rect 1140 -760 1180 -620
rect 1180 -760 1220 -620
rect 1220 -760 1230 -620
rect -190 -770 1230 -760
<< metal2 >>
rect -140 1370 1100 1390
rect -140 1210 -120 1370
rect 1090 1210 1100 1370
rect -140 960 1100 1210
rect -140 950 1090 960
rect -140 790 90 950
rect 150 790 510 950
rect 570 790 880 950
rect 940 790 1090 950
rect -140 780 1090 790
rect -230 480 1240 510
rect -230 320 10 480
rect 70 320 530 480
rect 590 320 1240 480
rect -230 -150 1240 320
rect -230 -310 400 -150
rect 460 -310 1240 -150
rect -230 -590 1240 -310
rect -230 -610 1250 -590
rect -230 -770 -190 -610
rect 1230 -770 1250 -610
rect -230 -790 1250 -770
<< labels >>
rlabel poly -270 200 -270 200 7 AIn
port 1 w
rlabel poly -270 -90 -270 -90 7 RST
port 2 w
rlabel space -510 -1289 -510 -1289 2 erase
rlabel poly 1290 -510 1290 -510 3 ENAD
port 3 e
rlabel poly 1290 120 1290 120 3 C+
port 4 e
rlabel poly 1280 720 1280 720 3 ENADb
port 5 e
rlabel locali 1280 1140 1280 1140 3 CompOut
port 6 e
rlabel poly -270 540 -270 540 7 Vb
port 7 w
<< end >>
