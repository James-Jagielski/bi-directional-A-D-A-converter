magic
tech sky130A
magscale 1 2
timestamp 1702611537
<< nwell >>
rect -760 90 -180 1260
rect -761 -469 -177 90
rect 4040 53 4620 1260
rect -760 -1875 -180 -469
rect 4038 -506 4622 53
rect 4040 -1905 4620 -506
<< nmos >>
rect 0 0 100 1200
rect 200 0 300 1200
rect 400 0 500 1200
rect 600 0 700 1200
rect 800 0 900 1200
rect 1000 0 1100 1200
rect 1200 0 1300 1200
rect 1400 0 1500 1200
rect 1770 0 1870 1200
rect 1970 0 2070 1200
rect 2340 0 2440 1200
rect 2540 0 2640 1200
rect 2740 0 2840 1200
rect 2940 0 3040 1200
rect 3140 0 3240 1200
rect 3340 0 3440 1200
rect 3540 0 3640 1200
rect 3740 0 3840 1200
rect 0 -1665 100 -465
rect 200 -1665 300 -465
rect 400 -1665 500 -465
rect 600 -1665 700 -465
rect 800 -1665 900 -465
rect 1000 -1665 1100 -465
rect 1200 -1665 1300 -465
rect 1400 -1665 1500 -465
rect 1770 -1665 1870 -465
rect 1970 -1665 2070 -465
rect 2340 -1665 2440 -465
rect 2540 -1665 2640 -465
rect 2740 -1665 2840 -465
rect 2940 -1665 3040 -465
rect 3140 -1665 3240 -465
rect 3340 -1665 3440 -465
rect 3540 -1665 3640 -465
rect 3740 -1665 3840 -465
<< pmos >>
rect -620 0 -520 1200
rect -420 0 -320 1200
rect 4180 0 4280 1200
rect 4380 0 4480 1200
rect -620 -1665 -520 -465
rect -420 -1665 -320 -465
rect 4180 -1665 4280 -465
rect 4380 -1665 4480 -465
<< ndiff >>
rect -100 1170 0 1200
rect -100 30 -70 1170
rect -30 30 0 1170
rect -100 0 0 30
rect 100 1170 200 1200
rect 100 30 130 1170
rect 170 30 200 1170
rect 100 0 200 30
rect 300 1170 400 1200
rect 300 30 330 1170
rect 370 30 400 1170
rect 300 0 400 30
rect 500 1170 600 1200
rect 500 30 530 1170
rect 570 30 600 1170
rect 500 0 600 30
rect 700 1170 800 1200
rect 700 30 730 1170
rect 770 30 800 1170
rect 700 0 800 30
rect 900 1170 1000 1200
rect 900 30 930 1170
rect 970 30 1000 1170
rect 900 0 1000 30
rect 1100 1170 1200 1200
rect 1100 30 1130 1170
rect 1170 30 1200 1170
rect 1100 0 1200 30
rect 1300 1170 1400 1200
rect 1300 30 1330 1170
rect 1370 30 1400 1170
rect 1300 0 1400 30
rect 1500 1170 1600 1200
rect 1500 30 1530 1170
rect 1570 30 1600 1170
rect 1500 0 1600 30
rect 1670 1170 1770 1200
rect 1670 30 1700 1170
rect 1740 30 1770 1170
rect 1670 0 1770 30
rect 1870 1170 1970 1200
rect 1870 30 1900 1170
rect 1940 30 1970 1170
rect 1870 0 1970 30
rect 2070 1170 2170 1200
rect 2070 30 2100 1170
rect 2140 30 2170 1170
rect 2070 0 2170 30
rect 2240 1170 2340 1200
rect 2240 30 2270 1170
rect 2310 30 2340 1170
rect 2240 0 2340 30
rect 2440 1170 2540 1200
rect 2440 30 2470 1170
rect 2510 30 2540 1170
rect 2440 0 2540 30
rect 2640 1170 2740 1200
rect 2640 30 2670 1170
rect 2710 30 2740 1170
rect 2640 0 2740 30
rect 2840 1170 2940 1200
rect 2840 30 2870 1170
rect 2910 30 2940 1170
rect 2840 0 2940 30
rect 3040 1170 3140 1200
rect 3040 30 3070 1170
rect 3110 30 3140 1170
rect 3040 0 3140 30
rect 3240 1170 3340 1200
rect 3240 30 3270 1170
rect 3310 30 3340 1170
rect 3240 0 3340 30
rect 3440 1170 3540 1200
rect 3440 30 3470 1170
rect 3510 30 3540 1170
rect 3440 0 3540 30
rect 3640 1170 3740 1200
rect 3640 30 3670 1170
rect 3710 30 3740 1170
rect 3640 0 3740 30
rect 3840 1170 3940 1200
rect 3840 30 3870 1170
rect 3910 30 3940 1170
rect 3840 0 3940 30
rect -100 -495 0 -465
rect -100 -1635 -70 -495
rect -30 -1635 0 -495
rect -100 -1665 0 -1635
rect 100 -495 200 -465
rect 100 -1635 130 -495
rect 170 -1635 200 -495
rect 100 -1665 200 -1635
rect 300 -495 400 -465
rect 300 -1635 330 -495
rect 370 -1635 400 -495
rect 300 -1665 400 -1635
rect 500 -495 600 -465
rect 500 -1635 530 -495
rect 570 -1635 600 -495
rect 500 -1665 600 -1635
rect 700 -495 800 -465
rect 700 -1635 730 -495
rect 770 -1635 800 -495
rect 700 -1665 800 -1635
rect 900 -495 1000 -465
rect 900 -1635 930 -495
rect 970 -1635 1000 -495
rect 900 -1665 1000 -1635
rect 1100 -495 1200 -465
rect 1100 -1635 1130 -495
rect 1170 -1635 1200 -495
rect 1100 -1665 1200 -1635
rect 1300 -495 1400 -465
rect 1300 -1635 1330 -495
rect 1370 -1635 1400 -495
rect 1300 -1665 1400 -1635
rect 1500 -495 1600 -465
rect 1500 -1635 1530 -495
rect 1570 -1635 1600 -495
rect 1500 -1665 1600 -1635
rect 1670 -495 1770 -465
rect 1670 -1635 1700 -495
rect 1740 -1635 1770 -495
rect 1670 -1665 1770 -1635
rect 1870 -495 1970 -465
rect 1870 -1635 1900 -495
rect 1940 -1635 1970 -495
rect 1870 -1665 1970 -1635
rect 2070 -495 2170 -465
rect 2070 -1635 2100 -495
rect 2140 -1635 2170 -495
rect 2070 -1665 2170 -1635
rect 2240 -495 2340 -465
rect 2240 -1635 2270 -495
rect 2310 -1635 2340 -495
rect 2240 -1665 2340 -1635
rect 2440 -495 2540 -465
rect 2440 -1635 2470 -495
rect 2510 -1635 2540 -495
rect 2440 -1665 2540 -1635
rect 2640 -495 2740 -465
rect 2640 -1635 2670 -495
rect 2710 -1635 2740 -495
rect 2640 -1665 2740 -1635
rect 2840 -495 2940 -465
rect 2840 -1635 2870 -495
rect 2910 -1635 2940 -495
rect 2840 -1665 2940 -1635
rect 3040 -495 3140 -465
rect 3040 -1635 3070 -495
rect 3110 -1635 3140 -495
rect 3040 -1665 3140 -1635
rect 3240 -495 3340 -465
rect 3240 -1635 3270 -495
rect 3310 -1635 3340 -495
rect 3240 -1665 3340 -1635
rect 3440 -495 3540 -465
rect 3440 -1635 3470 -495
rect 3510 -1635 3540 -495
rect 3440 -1665 3540 -1635
rect 3640 -495 3740 -465
rect 3640 -1635 3670 -495
rect 3710 -1635 3740 -495
rect 3640 -1665 3740 -1635
rect 3840 -495 3940 -465
rect 3840 -1635 3870 -495
rect 3910 -1635 3940 -495
rect 3840 -1665 3940 -1635
<< pdiff >>
rect -720 1170 -620 1200
rect -720 30 -690 1170
rect -650 30 -620 1170
rect -720 0 -620 30
rect -520 1170 -420 1200
rect -520 30 -490 1170
rect -450 30 -420 1170
rect -520 0 -420 30
rect -320 1170 -220 1200
rect -320 30 -290 1170
rect -250 30 -220 1170
rect -320 0 -220 30
rect 4080 1170 4180 1200
rect 4080 30 4110 1170
rect 4150 30 4180 1170
rect 4080 0 4180 30
rect 4280 1170 4380 1200
rect 4280 30 4310 1170
rect 4350 30 4380 1170
rect 4280 0 4380 30
rect 4480 1170 4580 1200
rect 4480 30 4510 1170
rect 4550 30 4580 1170
rect 4480 0 4580 30
rect -720 -495 -620 -465
rect -720 -1635 -690 -495
rect -650 -1635 -620 -495
rect -720 -1665 -620 -1635
rect -520 -495 -420 -465
rect -520 -1635 -490 -495
rect -450 -1635 -420 -495
rect -520 -1665 -420 -1635
rect -320 -495 -220 -465
rect -320 -1635 -290 -495
rect -250 -1635 -220 -495
rect -320 -1665 -220 -1635
rect 4080 -495 4180 -465
rect 4080 -1635 4110 -495
rect 4150 -1635 4180 -495
rect 4080 -1665 4180 -1635
rect 4280 -495 4380 -465
rect 4280 -1635 4310 -495
rect 4350 -1635 4380 -495
rect 4280 -1665 4380 -1635
rect 4480 -495 4580 -465
rect 4480 -1635 4510 -495
rect 4550 -1635 4580 -495
rect 4480 -1665 4580 -1635
<< ndiffc >>
rect -70 30 -30 1170
rect 130 30 170 1170
rect 330 30 370 1170
rect 530 30 570 1170
rect 730 30 770 1170
rect 930 30 970 1170
rect 1130 30 1170 1170
rect 1330 30 1370 1170
rect 1530 30 1570 1170
rect 1700 30 1740 1170
rect 1900 30 1940 1170
rect 2100 30 2140 1170
rect 2270 30 2310 1170
rect 2470 30 2510 1170
rect 2670 30 2710 1170
rect 2870 30 2910 1170
rect 3070 30 3110 1170
rect 3270 30 3310 1170
rect 3470 30 3510 1170
rect 3670 30 3710 1170
rect 3870 30 3910 1170
rect -70 -1635 -30 -495
rect 130 -1635 170 -495
rect 330 -1635 370 -495
rect 530 -1635 570 -495
rect 730 -1635 770 -495
rect 930 -1635 970 -495
rect 1130 -1635 1170 -495
rect 1330 -1635 1370 -495
rect 1530 -1635 1570 -495
rect 1700 -1635 1740 -495
rect 1900 -1635 1940 -495
rect 2100 -1635 2140 -495
rect 2270 -1635 2310 -495
rect 2470 -1635 2510 -495
rect 2670 -1635 2710 -495
rect 2870 -1635 2910 -495
rect 3070 -1635 3110 -495
rect 3270 -1635 3310 -495
rect 3470 -1635 3510 -495
rect 3670 -1635 3710 -495
rect 3870 -1635 3910 -495
<< pdiffc >>
rect -690 30 -650 1170
rect -490 30 -450 1170
rect -290 30 -250 1170
rect 4110 30 4150 1170
rect 4310 30 4350 1170
rect 4510 30 4550 1170
rect -690 -1635 -650 -495
rect -490 -1635 -450 -495
rect -290 -1635 -250 -495
rect 4110 -1635 4150 -495
rect 4310 -1635 4350 -495
rect 4510 -1635 4550 -495
<< psubdiff >>
rect 1840 -200 1980 -190
rect 1840 -240 1870 -200
rect 1950 -240 1980 -200
rect 1840 -250 1980 -240
rect 2099 -199 2241 -190
rect 2099 -239 2131 -199
rect 2211 -239 2241 -199
rect 2099 -250 2241 -239
rect 1266 -1844 1406 -1834
rect 1266 -1884 1296 -1844
rect 1376 -1884 1406 -1844
rect 1266 -1894 1406 -1884
<< nsubdiff >>
rect -530 -120 -390 -110
rect -530 -160 -500 -120
rect -420 -160 -390 -120
rect -530 -170 -390 -160
rect 4270 -150 4410 -140
rect 4270 -190 4300 -150
rect 4380 -190 4410 -150
rect 4270 -200 4410 -190
rect -530 -1785 -390 -1775
rect -530 -1825 -500 -1785
rect -420 -1825 -390 -1785
rect -530 -1835 -390 -1825
rect 4270 -1815 4410 -1805
rect 4270 -1855 4300 -1815
rect 4380 -1855 4410 -1815
rect 4270 -1865 4410 -1855
<< psubdiffcont >>
rect 1870 -240 1950 -200
rect 2131 -239 2211 -199
rect 1296 -1884 1376 -1844
<< nsubdiffcont >>
rect -500 -160 -420 -120
rect 4300 -190 4380 -150
rect -500 -1825 -420 -1785
rect 4300 -1855 4380 -1815
<< poly >>
rect -190 1290 -110 1310
rect -190 1250 -170 1290
rect -130 1280 -110 1290
rect 1880 1290 1960 1310
rect 1880 1280 1900 1290
rect -130 1250 1900 1280
rect 1940 1280 1960 1290
rect 3930 1290 4010 1300
rect 3930 1280 3950 1290
rect 1940 1250 3950 1280
rect 3990 1250 4010 1290
rect -620 1200 -520 1250
rect -420 1200 -320 1250
rect -190 1230 -110 1250
rect 0 1200 100 1250
rect 200 1200 300 1250
rect 400 1200 500 1250
rect 600 1200 700 1250
rect 800 1200 900 1250
rect 1000 1200 1100 1250
rect 1200 1200 1300 1250
rect 1400 1200 1500 1250
rect 1770 1230 2070 1250
rect 1770 1200 1870 1230
rect 1970 1200 2070 1230
rect 2340 1200 2440 1250
rect 2540 1200 2640 1250
rect 2740 1200 2840 1250
rect 2940 1200 3040 1250
rect 3140 1200 3240 1250
rect 3340 1200 3440 1250
rect 3540 1200 3640 1250
rect 3740 1200 3840 1250
rect 3930 1240 4010 1250
rect 4180 1200 4280 1250
rect 4380 1200 4480 1250
rect -620 -40 -520 0
rect -420 -30 -320 0
rect -420 -40 -50 -30
rect -620 -50 -50 -40
rect 0 -50 100 0
rect 200 -50 300 0
rect 400 -50 500 0
rect 600 -50 700 0
rect 800 -50 900 0
rect 1000 -50 1100 0
rect 1200 -50 1300 0
rect 1400 -50 1500 0
rect 1770 -50 1870 0
rect 1970 -50 2070 0
rect 2340 -50 2440 0
rect 2540 -50 2640 0
rect 2740 -50 2840 0
rect 2940 -50 3040 0
rect 3140 -50 3240 0
rect 3340 -50 3440 0
rect 3540 -50 3640 0
rect 3740 -50 3840 0
rect 4180 -30 4280 0
rect 4380 -30 4480 0
rect 3930 -50 4540 -30
rect -620 -70 -120 -50
rect -140 -100 -120 -70
rect -70 -100 -50 -50
rect -140 -120 -50 -100
rect 3930 -110 3950 -50
rect 4010 -70 4540 -50
rect 4010 -110 4030 -70
rect 3930 -130 4030 -110
rect -190 -375 -110 -355
rect -190 -415 -170 -375
rect -130 -385 -110 -375
rect 1880 -380 1960 -360
rect 1880 -385 1900 -380
rect -130 -415 1900 -385
rect -620 -465 -520 -415
rect -420 -465 -320 -415
rect -190 -435 -110 -415
rect 0 -465 100 -415
rect 200 -465 300 -415
rect 400 -465 500 -415
rect 600 -465 700 -415
rect 800 -465 900 -415
rect 1000 -465 1100 -415
rect 1200 -465 1300 -415
rect 1400 -465 1500 -415
rect 1770 -420 1900 -415
rect 1940 -385 1960 -380
rect 3930 -375 4010 -365
rect 3930 -385 3950 -375
rect 1940 -415 3950 -385
rect 3990 -415 4010 -375
rect 1940 -420 2070 -415
rect 1770 -440 2070 -420
rect 1770 -465 1870 -440
rect 1970 -465 2070 -440
rect 2340 -465 2440 -415
rect 2540 -465 2640 -415
rect 2740 -465 2840 -415
rect 2940 -465 3040 -415
rect 3140 -465 3240 -415
rect 3340 -465 3440 -415
rect 3540 -465 3640 -415
rect 3740 -465 3840 -415
rect 3930 -425 4010 -415
rect 4180 -465 4280 -415
rect 4380 -465 4480 -415
rect -620 -1705 -520 -1665
rect -420 -1695 -320 -1665
rect -420 -1705 -50 -1695
rect -620 -1715 -50 -1705
rect 0 -1715 100 -1665
rect 200 -1715 300 -1665
rect 400 -1715 500 -1665
rect 600 -1715 700 -1665
rect 800 -1715 900 -1665
rect 1000 -1715 1100 -1665
rect 1200 -1715 1300 -1665
rect 1400 -1715 1500 -1665
rect 1770 -1715 1870 -1665
rect 1970 -1715 2070 -1665
rect 2340 -1715 2440 -1665
rect 2540 -1715 2640 -1665
rect 2740 -1715 2840 -1665
rect 2940 -1715 3040 -1665
rect 3140 -1715 3240 -1665
rect 3340 -1715 3440 -1665
rect 3540 -1715 3640 -1665
rect 3740 -1715 3840 -1665
rect 3970 -1710 4080 -1690
rect 4180 -1705 4280 -1665
rect 4380 -1705 4480 -1665
rect 4180 -1710 4480 -1705
rect -620 -1735 -120 -1715
rect -140 -1765 -120 -1735
rect -70 -1765 -50 -1715
rect -140 -1785 -50 -1765
rect 3970 -1780 3990 -1710
rect 4060 -1750 4480 -1710
rect 4060 -1780 4080 -1750
rect 3970 -1800 4080 -1780
<< polycont >>
rect -170 1250 -130 1290
rect 1900 1250 1940 1290
rect 3950 1250 3990 1290
rect -120 -100 -70 -50
rect 3950 -110 4010 -50
rect -170 -415 -130 -375
rect 1900 -420 1940 -380
rect 3950 -415 3990 -375
rect -120 -1765 -70 -1715
rect 3990 -1780 4060 -1710
<< xpolycontact >>
rect 2339 -253 2779 -183
rect 2856 -253 3296 -183
rect 40 -1921 480 -1851
rect 564 -1921 1004 -1851
rect 1640 -1921 2080 -1851
rect 2164 -1921 2604 -1851
rect 2690 -1921 3130 -1851
rect 3214 -1921 3654 -1851
<< xpolyres >>
rect 2779 -253 2856 -183
rect 480 -1921 564 -1851
rect 2080 -1921 2164 -1851
rect 3130 -1921 3214 -1851
<< locali >>
rect -190 1290 -110 1310
rect -190 1280 -170 1290
rect -760 1250 -170 1280
rect -130 1250 -110 1290
rect -760 1230 -110 1250
rect 1880 1290 1960 1310
rect 1880 1250 1900 1290
rect 1940 1250 1960 1290
rect -270 1190 -230 1230
rect -710 1170 -630 1190
rect -710 30 -690 1170
rect -650 30 -630 1170
rect -710 10 -630 30
rect -510 1170 -430 1190
rect -510 30 -490 1170
rect -450 30 -430 1170
rect -510 10 -430 30
rect -310 1170 -230 1190
rect -310 30 -290 1170
rect -250 30 -230 1170
rect -310 10 -230 30
rect -90 1170 -10 1190
rect -90 30 -70 1170
rect -30 30 -10 1170
rect -90 10 -10 30
rect 110 1170 190 1190
rect 110 30 130 1170
rect 170 30 190 1170
rect 110 10 190 30
rect 310 1170 390 1190
rect 310 30 330 1170
rect 370 30 390 1170
rect 310 10 390 30
rect 510 1170 590 1190
rect 510 30 530 1170
rect 570 30 590 1170
rect 510 10 590 30
rect 710 1170 790 1190
rect 710 30 730 1170
rect 770 30 790 1170
rect 710 10 790 30
rect 910 1170 990 1190
rect 910 30 930 1170
rect 970 30 990 1170
rect 910 10 990 30
rect 1110 1170 1190 1190
rect 1110 30 1130 1170
rect 1170 30 1190 1170
rect 1110 10 1190 30
rect 1310 1170 1390 1190
rect 1310 30 1330 1170
rect 1370 30 1390 1170
rect 1310 10 1390 30
rect 1510 1170 1590 1190
rect 1510 30 1530 1170
rect 1570 30 1590 1170
rect 1510 10 1590 30
rect 1680 1170 1760 1190
rect 1680 30 1700 1170
rect 1740 30 1760 1170
rect 1680 10 1760 30
rect 1880 1170 1960 1250
rect 3930 1290 4010 1300
rect 3930 1250 3950 1290
rect 3990 1250 4130 1290
rect 3930 1240 4010 1250
rect 4090 1190 4130 1250
rect 1880 30 1900 1170
rect 1940 30 1960 1170
rect 1880 10 1960 30
rect 2080 1170 2160 1190
rect 2080 30 2100 1170
rect 2140 30 2160 1170
rect 2080 10 2160 30
rect 2250 1170 2330 1190
rect 2250 30 2270 1170
rect 2310 30 2330 1170
rect 2250 10 2330 30
rect 2450 1170 2530 1190
rect 2450 30 2470 1170
rect 2510 30 2530 1170
rect 2450 10 2530 30
rect 2650 1170 2730 1190
rect 2650 30 2670 1170
rect 2710 30 2730 1170
rect 2650 10 2730 30
rect 2850 1170 2930 1190
rect 2850 30 2870 1170
rect 2910 30 2930 1170
rect 2850 10 2930 30
rect 3050 1170 3130 1190
rect 3050 30 3070 1170
rect 3110 30 3130 1170
rect 3050 10 3130 30
rect 3250 1170 3330 1190
rect 3250 30 3270 1170
rect 3310 30 3330 1170
rect 3250 10 3330 30
rect 3450 1170 3530 1190
rect 3450 30 3470 1170
rect 3510 30 3530 1170
rect 3450 10 3530 30
rect 3650 1170 3730 1190
rect 3650 30 3670 1170
rect 3710 30 3730 1170
rect 3650 10 3730 30
rect 3850 1170 3930 1190
rect 3850 30 3870 1170
rect 3910 30 3930 1170
rect 3850 10 3930 30
rect 4090 1170 4170 1190
rect 4090 30 4110 1170
rect 4150 30 4170 1170
rect 4090 20 4170 30
rect 4290 1170 4370 1190
rect 4290 30 4310 1170
rect 4350 30 4370 1170
rect 4290 20 4370 30
rect 4490 1170 4570 1190
rect 4490 30 4510 1170
rect 4550 30 4570 1170
rect 4490 20 4570 30
rect -680 -30 -630 10
rect -60 -30 -10 10
rect 340 -30 390 10
rect 740 -30 790 10
rect 1140 -30 1190 10
rect 1540 -30 1590 10
rect 2280 -30 2330 10
rect 2680 -30 2730 10
rect 3080 -30 3130 10
rect 3480 -30 3530 10
rect 3880 -30 3930 10
rect 4490 -30 4540 20
rect -680 -50 4540 -30
rect -680 -70 -120 -50
rect -140 -100 -120 -70
rect -70 -80 3950 -50
rect -70 -100 -50 -80
rect -520 -120 -400 -110
rect -140 -120 -50 -100
rect 3930 -110 3950 -80
rect 4010 -80 4540 -50
rect 4010 -110 4030 -80
rect -520 -160 -500 -120
rect -420 -160 -400 -120
rect 3930 -130 4030 -110
rect -520 -170 -400 -160
rect 4280 -150 4400 -140
rect 1850 -200 1970 -190
rect 1850 -240 1870 -200
rect 1950 -240 1970 -200
rect 1850 -250 1970 -240
rect 2110 -199 2231 -190
rect 2110 -239 2131 -199
rect 2211 -239 2231 -199
rect 2110 -250 2231 -239
rect 4280 -190 4300 -150
rect 4380 -190 4400 -150
rect 4280 -200 4400 -190
rect -190 -375 -110 -355
rect -190 -395 -170 -375
rect -270 -400 -170 -395
rect -770 -415 -170 -400
rect -130 -415 -110 -375
rect -770 -435 -110 -415
rect 1880 -380 1960 -360
rect 1880 -420 1900 -380
rect 1940 -420 1960 -380
rect -770 -440 -230 -435
rect -270 -475 -230 -440
rect -710 -495 -630 -475
rect -710 -1635 -690 -495
rect -650 -1635 -630 -495
rect -710 -1655 -630 -1635
rect -510 -495 -430 -475
rect -510 -1635 -490 -495
rect -450 -1635 -430 -495
rect -510 -1655 -430 -1635
rect -310 -495 -230 -475
rect -310 -1635 -290 -495
rect -250 -1635 -230 -495
rect -310 -1655 -230 -1635
rect -90 -495 -10 -475
rect -90 -1635 -70 -495
rect -30 -1635 -10 -495
rect -90 -1655 -10 -1635
rect 110 -495 190 -475
rect 110 -1635 130 -495
rect 170 -1635 190 -495
rect 110 -1655 190 -1635
rect 310 -495 390 -475
rect 310 -1635 330 -495
rect 370 -1635 390 -495
rect 310 -1655 390 -1635
rect 510 -495 590 -475
rect 510 -1635 530 -495
rect 570 -1635 590 -495
rect 510 -1655 590 -1635
rect 710 -495 790 -475
rect 710 -1635 730 -495
rect 770 -1635 790 -495
rect 710 -1655 790 -1635
rect 910 -495 990 -475
rect 910 -1635 930 -495
rect 970 -1635 990 -495
rect 910 -1655 990 -1635
rect 1110 -495 1190 -475
rect 1110 -1635 1130 -495
rect 1170 -1635 1190 -495
rect 1110 -1655 1190 -1635
rect 1310 -495 1390 -475
rect 1310 -1635 1330 -495
rect 1370 -1635 1390 -495
rect 1310 -1655 1390 -1635
rect 1510 -495 1590 -475
rect 1510 -1635 1530 -495
rect 1570 -1635 1590 -495
rect 1510 -1655 1590 -1635
rect 1680 -495 1760 -475
rect 1680 -1635 1700 -495
rect 1740 -1635 1760 -495
rect 1680 -1655 1760 -1635
rect 1880 -495 1960 -420
rect 3930 -375 4010 -365
rect 3930 -415 3950 -375
rect 3990 -415 4130 -375
rect 3930 -425 4010 -415
rect 4090 -475 4130 -415
rect 1880 -1635 1900 -495
rect 1940 -1635 1960 -495
rect 1880 -1655 1960 -1635
rect 2080 -495 2160 -475
rect 2080 -1635 2100 -495
rect 2140 -1635 2160 -495
rect 2080 -1655 2160 -1635
rect 2250 -495 2330 -475
rect 2250 -1635 2270 -495
rect 2310 -1635 2330 -495
rect 2250 -1655 2330 -1635
rect 2450 -495 2530 -475
rect 2450 -1635 2470 -495
rect 2510 -1635 2530 -495
rect 2450 -1655 2530 -1635
rect 2650 -495 2730 -475
rect 2650 -1635 2670 -495
rect 2710 -1635 2730 -495
rect 2650 -1655 2730 -1635
rect 2850 -495 2930 -475
rect 2850 -1635 2870 -495
rect 2910 -1635 2930 -495
rect 2850 -1655 2930 -1635
rect 3050 -495 3130 -475
rect 3050 -1635 3070 -495
rect 3110 -1635 3130 -495
rect 3050 -1655 3130 -1635
rect 3250 -495 3330 -475
rect 3250 -1635 3270 -495
rect 3310 -1635 3330 -495
rect 3250 -1655 3330 -1635
rect 3450 -495 3530 -475
rect 3450 -1635 3470 -495
rect 3510 -1635 3530 -495
rect 3450 -1655 3530 -1635
rect 3650 -495 3730 -475
rect 3650 -1635 3670 -495
rect 3710 -1635 3730 -495
rect 3650 -1655 3730 -1635
rect 3850 -495 3930 -475
rect 3850 -1635 3870 -495
rect 3910 -1635 3930 -495
rect 3850 -1655 3930 -1635
rect 4090 -495 4170 -475
rect 4090 -1635 4110 -495
rect 4150 -1635 4170 -495
rect 4090 -1645 4170 -1635
rect 4290 -495 4370 -475
rect 4290 -1635 4310 -495
rect 4350 -1635 4370 -495
rect 4290 -1645 4370 -1635
rect 4490 -495 4570 -475
rect 4490 -1635 4510 -495
rect 4550 -1635 4570 -495
rect 4490 -1645 4570 -1635
rect -680 -1695 -630 -1655
rect -60 -1695 -10 -1655
rect 340 -1695 390 -1655
rect 740 -1695 790 -1655
rect 1140 -1695 1190 -1655
rect 1540 -1695 1590 -1655
rect 2280 -1695 2330 -1655
rect 2680 -1695 2730 -1655
rect 3080 -1695 3130 -1655
rect 3480 -1695 3530 -1655
rect 3880 -1695 3930 -1655
rect 3970 -1695 4080 -1690
rect 4490 -1695 4540 -1645
rect -680 -1710 4540 -1695
rect -680 -1715 3990 -1710
rect -680 -1735 -120 -1715
rect -140 -1765 -120 -1735
rect -70 -1745 3990 -1715
rect -70 -1765 -50 -1745
rect -520 -1785 -400 -1775
rect -140 -1785 -50 -1765
rect 3970 -1780 3990 -1745
rect 4060 -1745 4540 -1710
rect 4060 -1780 4080 -1745
rect -520 -1825 -500 -1785
rect -420 -1825 -400 -1785
rect 3970 -1800 4080 -1780
rect -520 -1835 -400 -1825
rect 4280 -1815 4400 -1805
rect 1276 -1844 1396 -1834
rect 1276 -1884 1296 -1844
rect 1376 -1884 1396 -1844
rect 1276 -1894 1396 -1884
rect 4280 -1855 4300 -1815
rect 4380 -1855 4400 -1815
rect 4280 -1865 4400 -1855
<< viali >>
rect -490 30 -450 1170
rect 130 30 170 1170
rect 530 30 570 1170
rect 930 30 970 1170
rect 1330 30 1370 1170
rect 1700 30 1740 1170
rect 2100 30 2140 1170
rect 2470 30 2510 1170
rect 2870 30 2910 1170
rect 3270 30 3310 1170
rect 3670 30 3710 1170
rect 4310 30 4350 1170
rect -500 -160 -420 -120
rect 1870 -240 1950 -200
rect 2131 -239 2211 -199
rect 2339 -253 2779 -183
rect 2856 -253 3296 -183
rect 4300 -190 4380 -150
rect -490 -1635 -450 -495
rect 130 -1635 170 -495
rect 530 -1635 570 -495
rect 930 -1635 970 -495
rect 1330 -1635 1370 -495
rect 1700 -1635 1740 -495
rect 2100 -1635 2140 -495
rect 2470 -1635 2510 -495
rect 2870 -1635 2910 -495
rect 3270 -1635 3310 -495
rect 3670 -1635 3710 -495
rect 4310 -1635 4350 -495
rect -500 -1825 -420 -1785
rect 40 -1921 480 -1851
rect 564 -1921 1004 -1851
rect 1296 -1884 1376 -1844
rect 1640 -1921 2080 -1851
rect 2164 -1921 2604 -1851
rect 2690 -1921 3130 -1851
rect 3214 -1921 3654 -1851
rect 4300 -1855 4380 -1815
<< metal1 >>
rect -510 1180 -430 1190
rect -510 20 -500 1180
rect -440 20 -430 1180
rect -510 10 -430 20
rect -100 1170 1600 1200
rect -100 30 130 1170
rect 170 30 530 1170
rect 570 30 930 1170
rect 970 30 1330 1170
rect 1370 30 1600 1170
rect -100 0 1600 30
rect 1670 1190 2170 1200
rect 1670 10 1680 1190
rect 1760 10 2080 1190
rect 2160 10 2170 1190
rect 1670 0 2170 10
rect 2240 1170 3940 1200
rect 2240 30 2470 1170
rect 2510 30 2870 1170
rect 2910 30 3270 1170
rect 3310 30 3670 1170
rect 3710 30 3940 1170
rect 2240 0 3940 30
rect 4290 1180 4370 1190
rect 4290 20 4300 1180
rect 4360 20 4370 1180
rect 4290 10 4370 20
rect 1510 -60 1600 0
rect 2250 -60 2330 0
rect 1510 -100 2330 -60
rect -530 -160 -500 -100
rect -420 -160 -390 -100
rect -530 -170 -390 -160
rect 3240 -163 3317 0
rect 2326 -183 2799 -163
rect 1840 -250 1850 -190
rect 1970 -250 1980 -190
rect 2099 -250 2110 -190
rect 2231 -250 2241 -190
rect 2326 -253 2339 -183
rect 2779 -253 2799 -183
rect 2326 -265 2799 -253
rect 2846 -164 3317 -163
rect 2846 -183 3316 -164
rect 2846 -253 2856 -183
rect 3296 -253 3316 -183
rect 4270 -200 4280 -130
rect 4380 -200 4410 -130
rect 2327 -266 2782 -265
rect 2846 -266 3316 -253
rect 2520 -465 2603 -454
rect -510 -485 -430 -475
rect -510 -1645 -500 -485
rect -440 -1645 -430 -485
rect -510 -1655 -430 -1645
rect -100 -495 1600 -465
rect -100 -1635 130 -495
rect 170 -1635 530 -495
rect 570 -1635 930 -495
rect 970 -1635 1330 -495
rect 1370 -1635 1600 -495
rect -100 -1665 1600 -1635
rect 1670 -475 2170 -465
rect 1670 -1655 1680 -475
rect 1760 -1655 2080 -475
rect 2160 -1655 2170 -475
rect 1670 -1660 2170 -1655
rect 2240 -495 3940 -465
rect 2240 -1635 2470 -495
rect 2510 -1635 2870 -495
rect 2910 -1635 3270 -495
rect 3310 -1635 3670 -495
rect 3710 -1635 3940 -495
rect 2240 -1660 3940 -1635
rect 4290 -485 4370 -475
rect 4290 -1645 4300 -485
rect 4360 -1645 4370 -485
rect 4290 -1655 4370 -1645
rect 928 -1710 1012 -1665
rect -530 -1825 -500 -1765
rect -420 -1825 -390 -1765
rect -530 -1835 -390 -1825
rect 928 -1833 1010 -1710
rect 1510 -1730 1600 -1665
rect 2250 -1665 3940 -1660
rect 2250 -1730 2330 -1665
rect 1510 -1796 2330 -1730
rect 1510 -1797 1863 -1796
rect 2036 -1797 2330 -1796
rect 2520 -1745 2616 -1665
rect 2520 -1829 2615 -1745
rect 406 -1838 494 -1837
rect 28 -1851 494 -1838
rect 28 -1921 40 -1851
rect 480 -1921 494 -1851
rect 28 -1934 494 -1921
rect 406 -1935 494 -1934
rect 552 -1840 1010 -1833
rect 552 -1851 1012 -1840
rect 552 -1921 564 -1851
rect 1004 -1921 1012 -1851
rect 1260 -1890 1270 -1830
rect 1400 -1890 1410 -1830
rect 1869 -1837 1971 -1836
rect 1869 -1838 2092 -1837
rect 1260 -1891 1276 -1890
rect 1394 -1891 1410 -1890
rect 1260 -1900 1410 -1891
rect 1628 -1851 2092 -1838
rect 552 -1940 1012 -1921
rect 1628 -1921 1640 -1851
rect 2080 -1921 2092 -1851
rect 1628 -1934 2092 -1921
rect 1930 -1936 2092 -1934
rect 2156 -1851 2615 -1829
rect 3202 -1830 3286 -1665
rect 3202 -1831 3664 -1830
rect 2156 -1921 2164 -1851
rect 2604 -1921 2615 -1851
rect 2156 -1938 2615 -1921
rect 2678 -1851 3142 -1839
rect 2678 -1921 2690 -1851
rect 3130 -1921 3142 -1851
rect 2678 -1934 3142 -1921
rect 3203 -1851 3664 -1831
rect 3203 -1921 3214 -1851
rect 3654 -1921 3664 -1851
rect 4270 -1855 4300 -1795
rect 4380 -1855 4410 -1795
rect 4270 -1865 4410 -1855
rect 3203 -1937 3664 -1921
<< via1 >>
rect -500 1170 -440 1180
rect -500 30 -490 1170
rect -490 30 -450 1170
rect -450 30 -440 1170
rect -500 20 -440 30
rect 1680 1170 1760 1190
rect 1680 30 1700 1170
rect 1700 30 1740 1170
rect 1740 30 1760 1170
rect 1680 10 1760 30
rect 2080 1170 2160 1190
rect 2080 30 2100 1170
rect 2100 30 2140 1170
rect 2140 30 2160 1170
rect 2080 10 2160 30
rect 4300 1170 4360 1180
rect 4300 30 4310 1170
rect 4310 30 4350 1170
rect 4350 30 4360 1170
rect 4300 20 4360 30
rect -500 -120 -420 -100
rect -500 -160 -420 -120
rect 1850 -200 1970 -190
rect 1850 -240 1870 -200
rect 1870 -240 1950 -200
rect 1950 -240 1970 -200
rect 1850 -250 1970 -240
rect 2110 -199 2231 -190
rect 2110 -239 2131 -199
rect 2131 -239 2211 -199
rect 2211 -239 2231 -199
rect 2110 -250 2231 -239
rect 2339 -253 2779 -183
rect 4280 -150 4380 -130
rect 4280 -190 4300 -150
rect 4300 -190 4380 -150
rect 4280 -200 4380 -190
rect -500 -495 -440 -485
rect -500 -1635 -490 -495
rect -490 -1635 -450 -495
rect -450 -1635 -440 -495
rect -500 -1645 -440 -1635
rect 1680 -495 1760 -475
rect 1680 -1635 1700 -495
rect 1700 -1635 1740 -495
rect 1740 -1635 1760 -495
rect 1680 -1655 1760 -1635
rect 2080 -495 2160 -475
rect 2080 -1635 2100 -495
rect 2100 -1635 2140 -495
rect 2140 -1635 2160 -495
rect 2080 -1655 2160 -1635
rect 4300 -495 4360 -485
rect 4300 -1635 4310 -495
rect 4310 -1635 4350 -495
rect 4350 -1635 4360 -495
rect 4300 -1645 4360 -1635
rect -500 -1785 -420 -1765
rect -500 -1825 -420 -1785
rect 40 -1921 480 -1851
rect 1270 -1844 1400 -1830
rect 1270 -1884 1296 -1844
rect 1296 -1884 1376 -1844
rect 1376 -1884 1400 -1844
rect 1270 -1890 1400 -1884
rect 1276 -1891 1394 -1890
rect 1640 -1921 2080 -1851
rect 2690 -1921 3130 -1851
rect 4300 -1815 4380 -1795
rect 4300 -1855 4380 -1815
<< metal2 >>
rect -760 1270 4380 1320
rect -520 1180 -420 1270
rect -520 20 -500 1180
rect -440 20 -420 1180
rect -520 -100 -420 20
rect 1670 1190 2170 1200
rect 1670 10 1680 1190
rect 1760 10 2080 1190
rect 2160 10 2170 1190
rect 1670 0 2170 10
rect 4280 1180 4380 1270
rect 4280 20 4300 1180
rect 4360 20 4380 1180
rect -520 -160 -500 -100
rect -420 -160 -400 -110
rect -520 -170 -400 -160
rect 1830 -163 1990 0
rect 4280 -130 4380 20
rect -520 -485 -420 -170
rect 1830 -183 2799 -163
rect 1830 -190 2339 -183
rect 1830 -250 1850 -190
rect 1970 -250 2110 -190
rect 2231 -250 2339 -190
rect 1830 -253 2339 -250
rect 2779 -253 2799 -183
rect 1830 -265 2799 -253
rect 4380 -200 4400 -140
rect 1830 -465 1990 -265
rect -520 -1645 -500 -485
rect -440 -1645 -420 -485
rect -520 -1765 -420 -1645
rect 1670 -475 2170 -465
rect 1670 -1655 1680 -475
rect 1760 -1655 2080 -475
rect 2160 -1655 2170 -475
rect 1670 -1665 2170 -1655
rect 4280 -485 4380 -200
rect 4280 -1645 4300 -485
rect 4360 -1645 4380 -485
rect 1830 -1666 1990 -1665
rect 1869 -1704 1971 -1666
rect 1870 -1748 1970 -1704
rect -520 -1825 -500 -1765
rect -420 -1825 -400 -1775
rect -520 -1835 -400 -1825
rect 406 -1807 2766 -1748
rect 406 -1837 494 -1807
rect 28 -1851 494 -1837
rect 28 -1880 40 -1851
rect -770 -1921 40 -1880
rect 480 -1921 494 -1851
rect 1260 -1830 1408 -1807
rect 1260 -1890 1270 -1830
rect 1400 -1890 1408 -1830
rect 1260 -1891 1276 -1890
rect 1394 -1891 1408 -1890
rect 1260 -1895 1408 -1891
rect 1628 -1851 2094 -1807
rect -770 -1935 494 -1921
rect 1628 -1921 1640 -1851
rect 2080 -1921 2094 -1851
rect 1628 -1935 2094 -1921
rect 2678 -1839 2766 -1807
rect 4280 -1795 4380 -1645
rect 2678 -1851 3143 -1839
rect 2678 -1921 2690 -1851
rect 3130 -1921 3143 -1851
rect 4280 -1855 4300 -1795
rect 4380 -1855 4400 -1805
rect 4280 -1865 4400 -1855
rect 2678 -1935 3143 -1921
rect -770 -1940 30 -1935
rect 1930 -1936 2094 -1935
<< labels >>
rlabel locali -760 1260 -760 1260 7 Vb
port 1 w
rlabel locali -770 -420 -770 -420 7 Vcp
port 2 w
rlabel metal2 -760 1300 -760 1300 7 VDD
port 3 w
rlabel metal2 -770 -1910 -770 -1910 7 GND
port 4 w
<< end >>
