magic
tech sky130A
timestamp 1702586952
<< nwell >>
rect -175 -20 780 120
<< nmos >>
rect -60 -190 -45 -90
rect 85 -190 100 -90
rect 150 -190 165 -90
rect 295 -190 310 -90
rect 440 -190 455 -90
rect 505 -190 520 -90
rect 650 -190 665 -90
rect -125 -385 -110 -285
rect -60 -385 -45 -285
rect 5 -385 20 -285
rect 195 -385 210 -285
rect 260 -385 275 -285
rect 330 -385 345 -285
rect 395 -385 410 -285
rect 585 -385 600 -285
rect 650 -385 665 -285
rect 715 -385 730 -285
<< pmos >>
rect -105 0 -90 100
rect -40 0 -25 100
rect 25 0 40 100
rect 90 0 105 100
rect 155 0 170 100
rect 220 0 235 100
rect 370 0 385 100
rect 435 0 450 100
rect 500 0 515 100
rect 565 0 580 100
rect 630 0 645 100
rect 695 0 710 100
<< ndiff >>
rect -110 -105 -60 -90
rect -110 -175 -95 -105
rect -75 -175 -60 -105
rect -110 -190 -60 -175
rect -45 -105 5 -90
rect -45 -175 -30 -105
rect -10 -175 5 -105
rect -45 -190 5 -175
rect 35 -105 85 -90
rect 35 -175 50 -105
rect 70 -175 85 -105
rect 35 -190 85 -175
rect 100 -105 150 -90
rect 100 -175 115 -105
rect 135 -175 150 -105
rect 100 -190 150 -175
rect 165 -105 215 -90
rect 165 -175 180 -105
rect 200 -175 215 -105
rect 165 -190 215 -175
rect 245 -105 295 -90
rect 245 -175 260 -105
rect 280 -175 295 -105
rect 245 -190 295 -175
rect 310 -105 360 -90
rect 310 -175 325 -105
rect 345 -175 360 -105
rect 310 -190 360 -175
rect 390 -105 440 -90
rect 390 -175 405 -105
rect 425 -175 440 -105
rect 390 -190 440 -175
rect 455 -105 505 -90
rect 455 -175 470 -105
rect 490 -175 505 -105
rect 455 -190 505 -175
rect 520 -105 570 -90
rect 520 -175 535 -105
rect 555 -175 570 -105
rect 520 -190 570 -175
rect 600 -105 650 -90
rect 600 -175 615 -105
rect 635 -175 650 -105
rect 600 -190 650 -175
rect 665 -105 715 -90
rect 665 -175 680 -105
rect 700 -175 715 -105
rect 665 -190 715 -175
rect -175 -300 -125 -285
rect -175 -370 -160 -300
rect -140 -370 -125 -300
rect -175 -385 -125 -370
rect -110 -300 -60 -285
rect -110 -370 -95 -300
rect -75 -370 -60 -300
rect -110 -385 -60 -370
rect -45 -300 5 -285
rect -45 -370 -30 -300
rect -10 -370 5 -300
rect -45 -385 5 -370
rect 20 -300 70 -285
rect 20 -370 35 -300
rect 55 -370 70 -300
rect 20 -385 70 -370
rect 145 -300 195 -285
rect 145 -370 160 -300
rect 180 -370 195 -300
rect 145 -385 195 -370
rect 210 -300 260 -285
rect 210 -370 225 -300
rect 245 -370 260 -300
rect 210 -385 260 -370
rect 275 -300 330 -285
rect 275 -370 290 -300
rect 315 -370 330 -300
rect 275 -385 330 -370
rect 345 -300 395 -285
rect 345 -370 360 -300
rect 380 -370 395 -300
rect 345 -385 395 -370
rect 410 -300 460 -285
rect 410 -370 425 -300
rect 445 -370 460 -300
rect 410 -385 460 -370
rect 535 -300 585 -285
rect 535 -370 550 -300
rect 570 -370 585 -300
rect 535 -385 585 -370
rect 600 -300 650 -285
rect 600 -370 615 -300
rect 635 -370 650 -300
rect 600 -385 650 -370
rect 665 -300 715 -285
rect 665 -370 680 -300
rect 700 -370 715 -300
rect 665 -385 715 -370
rect 730 -300 780 -285
rect 730 -370 745 -300
rect 765 -370 780 -300
rect 730 -385 780 -370
<< pdiff >>
rect -155 85 -105 100
rect -155 15 -140 85
rect -120 15 -105 85
rect -155 0 -105 15
rect -90 85 -40 100
rect -90 15 -75 85
rect -55 15 -40 85
rect -90 0 -40 15
rect -25 85 25 100
rect -25 15 -10 85
rect 10 15 25 85
rect -25 0 25 15
rect 40 85 90 100
rect 40 15 55 85
rect 75 15 90 85
rect 40 0 90 15
rect 105 0 155 100
rect 170 85 220 100
rect 170 15 185 85
rect 205 15 220 85
rect 170 0 220 15
rect 235 85 285 100
rect 235 15 250 85
rect 270 15 285 85
rect 235 0 285 15
rect 320 85 370 100
rect 320 15 335 85
rect 355 15 370 85
rect 320 0 370 15
rect 385 85 435 100
rect 385 15 400 85
rect 420 15 435 85
rect 385 0 435 15
rect 450 0 500 100
rect 515 85 565 100
rect 515 15 530 85
rect 550 15 565 85
rect 515 0 565 15
rect 580 85 630 100
rect 580 15 595 85
rect 615 15 630 85
rect 580 0 630 15
rect 645 85 695 100
rect 645 15 660 85
rect 680 15 695 85
rect 645 0 695 15
rect 710 85 760 100
rect 710 15 725 85
rect 745 15 760 85
rect 710 0 760 15
<< ndiffc >>
rect -95 -175 -75 -105
rect -30 -175 -10 -105
rect 50 -175 70 -105
rect 115 -175 135 -105
rect 180 -175 200 -105
rect 260 -175 280 -105
rect 325 -175 345 -105
rect 405 -175 425 -105
rect 470 -175 490 -105
rect 535 -175 555 -105
rect 615 -175 635 -105
rect 680 -175 700 -105
rect -160 -370 -140 -300
rect -95 -370 -75 -300
rect -30 -370 -10 -300
rect 35 -370 55 -300
rect 160 -370 180 -300
rect 225 -370 245 -300
rect 290 -370 315 -300
rect 360 -370 380 -300
rect 425 -370 445 -300
rect 550 -370 570 -300
rect 615 -370 635 -300
rect 680 -370 700 -300
rect 745 -370 765 -300
<< pdiffc >>
rect -140 15 -120 85
rect -75 15 -55 85
rect -10 15 10 85
rect 55 15 75 85
rect 185 15 205 85
rect 250 15 270 85
rect 335 15 355 85
rect 400 15 420 85
rect 530 15 550 85
rect 595 15 615 85
rect 660 15 680 85
rect 725 15 745 85
<< poly >>
rect -105 100 -90 115
rect -40 100 -25 115
rect 25 100 40 115
rect 90 100 105 115
rect 155 100 170 115
rect 220 100 235 115
rect 370 100 385 115
rect 435 100 450 115
rect 500 100 515 115
rect 565 100 580 115
rect 630 100 645 115
rect 695 100 710 115
rect -105 -15 -90 0
rect -40 -15 -25 0
rect 25 -15 40 0
rect 90 -15 105 0
rect 155 -15 170 0
rect 220 -15 235 0
rect 370 -15 385 0
rect 435 -15 450 0
rect 500 -15 515 0
rect 565 -15 580 0
rect 630 -15 645 0
rect 695 -15 710 0
rect -60 -90 -45 -75
rect 85 -90 100 -75
rect 150 -90 165 -75
rect 295 -90 310 -70
rect 440 -90 455 -75
rect 505 -90 520 -75
rect 650 -90 665 -75
rect -60 -205 -45 -190
rect 85 -205 100 -190
rect 150 -200 165 -190
rect -85 -215 -45 -205
rect 150 -215 210 -200
rect 295 -205 310 -190
rect 440 -200 455 -190
rect -85 -235 -75 -215
rect -55 -235 -45 -215
rect -85 -245 -45 -235
rect -125 -285 -110 -270
rect -60 -285 -45 -270
rect 5 -285 20 -270
rect 195 -285 210 -215
rect 395 -215 455 -200
rect 505 -205 520 -190
rect 650 -205 665 -190
rect 650 -215 690 -205
rect 260 -285 275 -270
rect 330 -285 345 -270
rect 395 -285 410 -215
rect 650 -235 660 -215
rect 680 -235 690 -215
rect 650 -245 690 -235
rect 585 -285 600 -270
rect 650 -285 665 -270
rect 715 -285 730 -270
rect -125 -400 -110 -385
rect -60 -400 -45 -385
rect 5 -400 20 -385
rect 195 -425 210 -385
rect 260 -400 275 -385
rect 330 -400 345 -385
rect 395 -425 410 -385
rect 585 -400 600 -385
rect 650 -400 665 -385
rect 715 -400 730 -385
rect 195 -440 410 -425
<< polycont >>
rect -75 -235 -55 -215
rect 660 -235 680 -215
<< locali >>
rect -150 85 -110 95
rect -150 25 -140 85
rect -185 15 -140 25
rect -120 15 -110 85
rect -185 5 -110 15
rect -85 85 20 95
rect -85 15 -75 85
rect -55 15 -10 85
rect 10 15 20 85
rect -85 5 20 15
rect 45 85 85 95
rect 45 15 55 85
rect 75 15 85 85
rect 45 5 85 15
rect 175 85 215 95
rect 175 15 185 85
rect 205 15 215 85
rect 175 5 215 15
rect 240 85 280 95
rect 240 15 250 85
rect 270 15 280 85
rect 240 5 280 15
rect 325 85 365 95
rect 325 15 335 85
rect 355 15 365 85
rect 325 5 365 15
rect 390 85 430 95
rect 390 15 400 85
rect 420 15 430 85
rect 390 5 430 15
rect 520 85 560 95
rect 520 15 530 85
rect 550 15 560 85
rect 520 5 560 15
rect 585 85 690 95
rect 585 15 595 85
rect 615 15 660 85
rect 680 15 690 85
rect 585 5 690 15
rect 715 85 755 95
rect 715 15 725 85
rect 745 25 755 85
rect 745 15 790 25
rect 715 5 790 15
rect -185 -290 -165 5
rect -85 -15 -65 5
rect -145 -35 -65 -15
rect 670 -15 690 5
rect 670 -35 750 -15
rect -145 -205 -125 -35
rect -85 -75 -55 -55
rect -85 -95 -65 -75
rect -105 -105 -65 -95
rect -105 -175 -95 -105
rect -75 -175 -65 -105
rect -105 -185 -65 -175
rect -40 -105 0 -95
rect -40 -175 -30 -105
rect -10 -175 0 -105
rect -40 -185 0 -175
rect 40 -105 80 -95
rect 40 -175 50 -105
rect 70 -175 80 -105
rect 40 -185 80 -175
rect 105 -105 145 -95
rect 105 -175 115 -105
rect 135 -175 145 -105
rect 105 -185 145 -175
rect 170 -105 210 -95
rect 170 -175 180 -105
rect 200 -175 210 -105
rect 170 -185 210 -175
rect 250 -105 290 -95
rect 250 -175 260 -105
rect 280 -175 290 -105
rect 250 -185 290 -175
rect 315 -105 355 -95
rect 315 -175 325 -105
rect 345 -175 355 -105
rect 315 -185 355 -175
rect 395 -105 435 -95
rect 395 -175 405 -105
rect 425 -175 435 -105
rect 395 -185 435 -175
rect 460 -105 500 -95
rect 460 -175 470 -105
rect 490 -175 500 -105
rect 460 -185 500 -175
rect 525 -105 565 -95
rect 525 -175 535 -105
rect 555 -175 565 -105
rect 525 -185 565 -175
rect 605 -105 645 -95
rect 605 -175 615 -105
rect 635 -175 645 -105
rect 605 -185 645 -175
rect 670 -105 710 -95
rect 670 -175 680 -105
rect 700 -175 710 -105
rect 670 -185 710 -175
rect 730 -205 750 -35
rect -145 -215 -45 -205
rect -145 -225 -75 -215
rect -85 -235 -75 -225
rect -55 -235 -45 -215
rect -85 -245 -45 -235
rect 650 -215 750 -205
rect 650 -235 660 -215
rect 680 -225 750 -215
rect 680 -235 690 -225
rect 650 -245 690 -235
rect -85 -290 -65 -245
rect 670 -290 690 -245
rect 770 -290 790 5
rect -185 -300 -130 -290
rect -185 -310 -160 -300
rect -170 -370 -160 -310
rect -140 -370 -130 -300
rect -170 -380 -130 -370
rect -105 -300 0 -290
rect -105 -370 -95 -300
rect -75 -370 -30 -300
rect -10 -370 0 -300
rect -105 -380 0 -370
rect 25 -300 65 -290
rect 25 -370 35 -300
rect 55 -370 65 -300
rect 25 -380 65 -370
rect 150 -300 190 -290
rect 150 -370 160 -300
rect 180 -370 190 -300
rect 150 -380 190 -370
rect 215 -300 255 -290
rect 215 -370 225 -300
rect 245 -370 255 -300
rect 215 -380 255 -370
rect 280 -300 325 -290
rect 280 -370 290 -300
rect 315 -370 325 -300
rect 280 -380 325 -370
rect 350 -300 390 -290
rect 350 -370 360 -300
rect 380 -370 390 -300
rect 350 -380 390 -370
rect 415 -300 455 -290
rect 415 -370 425 -300
rect 445 -370 455 -300
rect 415 -380 455 -370
rect 540 -300 580 -290
rect 540 -370 550 -300
rect 570 -370 580 -300
rect 540 -380 580 -370
rect 605 -300 710 -290
rect 605 -370 615 -300
rect 635 -370 680 -300
rect 700 -370 710 -300
rect 605 -380 710 -370
rect 735 -300 790 -290
rect 735 -370 745 -300
rect 765 -310 790 -300
rect 765 -370 775 -310
rect 735 -380 775 -370
<< viali >>
rect 185 15 205 85
rect 400 15 420 85
rect 260 -175 280 -105
rect 160 -370 180 -300
rect 425 -370 445 -300
<< metal1 >>
rect 175 90 215 95
rect 175 10 180 90
rect 210 10 215 90
rect 175 5 215 10
rect 390 90 430 95
rect 390 10 395 90
rect 425 10 430 90
rect 390 5 430 10
rect 250 -100 290 -95
rect 250 -180 255 -100
rect 285 -180 290 -100
rect 250 -185 290 -180
rect 150 -295 190 -290
rect 150 -375 155 -295
rect 185 -375 190 -295
rect 150 -380 190 -375
rect 415 -295 455 -290
rect 415 -375 420 -295
rect 450 -375 455 -295
rect 415 -380 455 -375
<< via1 >>
rect 180 85 210 90
rect 180 15 185 85
rect 185 15 205 85
rect 205 15 210 85
rect 180 10 210 15
rect 395 85 425 90
rect 395 15 400 85
rect 400 15 420 85
rect 420 15 425 85
rect 395 10 425 15
rect 255 -105 285 -100
rect 255 -175 260 -105
rect 260 -175 280 -105
rect 280 -175 285 -105
rect 255 -180 285 -175
rect 155 -300 185 -295
rect 155 -370 160 -300
rect 160 -370 180 -300
rect 180 -370 185 -300
rect 155 -375 185 -370
rect 420 -300 450 -295
rect 420 -370 425 -300
rect 425 -370 445 -300
rect 445 -370 450 -300
rect 420 -375 450 -370
<< metal2 >>
rect 175 90 215 95
rect 175 10 180 90
rect 210 10 215 90
rect 175 5 215 10
rect 390 90 430 95
rect 390 10 395 90
rect 425 10 430 90
rect 390 5 430 10
rect 250 -100 290 -95
rect 250 -180 255 -100
rect 285 -180 290 -100
rect 250 -185 290 -180
rect 150 -295 190 -290
rect 150 -375 155 -295
rect 185 -375 190 -295
rect 150 -380 190 -375
rect 415 -295 455 -290
rect 415 -375 420 -295
rect 450 -375 455 -295
rect 415 -380 455 -375
<< end >>
