magic
tech sky130A
timestamp 1702595637
<< metal3 >>
rect 1685 880 6770 1015
rect 1685 -15 6715 880
rect 6615 -70 6770 -65
rect 1685 -205 6770 -70
rect 1685 -1100 6715 -205
rect 1685 -1295 6770 -1155
rect 1685 -2185 6715 -1295
rect 1685 -2380 6770 -2240
rect 1685 -3270 6715 -2380
rect 1685 -3455 6770 -3325
rect 1685 -3640 6770 -3510
rect 1685 -3825 6770 -3695
rect 1685 -4010 6770 -3880
rect 1685 -4195 6770 -4065
rect 1685 -4380 6770 -4250
<< mimcap >>
rect 1700 990 6700 1000
rect 1700 955 1710 990
rect 1745 955 6700 990
rect 1700 0 6700 955
rect 1700 -95 6700 -85
rect 1700 -130 1710 -95
rect 1745 -130 6700 -95
rect 1700 -1085 6700 -130
rect 1700 -1180 6700 -1170
rect 1700 -1215 1710 -1180
rect 1745 -1215 6700 -1180
rect 1700 -2170 6700 -1215
rect 1700 -2265 6700 -2255
rect 1700 -2300 1710 -2265
rect 1745 -2300 6700 -2265
rect 1700 -3255 6700 -2300
rect 1700 -3350 6700 -3340
rect 1700 -3385 1710 -3350
rect 1745 -3385 6700 -3350
rect 1700 -3440 6700 -3385
rect 1700 -3535 6700 -3525
rect 1700 -3570 1710 -3535
rect 1745 -3570 6700 -3535
rect 1700 -3625 6700 -3570
rect 1700 -3720 6700 -3710
rect 1700 -3755 1710 -3720
rect 1745 -3755 6700 -3720
rect 1700 -3810 6700 -3755
rect 1700 -3905 6700 -3895
rect 1700 -3940 1710 -3905
rect 1745 -3940 6700 -3905
rect 1700 -3995 6700 -3940
rect 1700 -4090 6700 -4080
rect 1700 -4125 1710 -4090
rect 1745 -4125 6700 -4090
rect 1700 -4180 6700 -4125
rect 1700 -4275 6700 -4265
rect 1700 -4310 1710 -4275
rect 1745 -4310 6700 -4275
rect 1700 -4365 6700 -4310
<< mimcapcontact >>
rect 1710 955 1745 990
rect 1710 -130 1745 -95
rect 1710 -1215 1745 -1180
rect 1710 -2300 1745 -2265
rect 1710 -3385 1745 -3350
rect 1710 -3570 1745 -3535
rect 1710 -3755 1745 -3720
rect 1710 -3940 1745 -3905
rect 1710 -4125 1745 -4090
rect 1710 -4310 1745 -4275
<< metal4 >>
rect 1630 990 1750 1000
rect 1630 955 1710 990
rect 1745 955 1750 990
rect 1630 950 1750 955
rect 1630 -95 1750 -85
rect 1630 -130 1710 -95
rect 1745 -130 1750 -95
rect 1630 -135 1750 -130
rect 1630 -1180 1750 -1170
rect 1630 -1215 1710 -1180
rect 1745 -1215 1750 -1180
rect 1630 -1220 1750 -1215
rect 1630 -2265 1750 -2255
rect 1630 -2300 1710 -2265
rect 1745 -2300 1750 -2265
rect 1630 -2305 1750 -2300
rect 1630 -3350 1750 -3340
rect 1630 -3385 1710 -3350
rect 1745 -3385 1750 -3350
rect 1630 -3390 1750 -3385
rect 1630 -3535 1750 -3525
rect 1630 -3570 1710 -3535
rect 1745 -3570 1750 -3535
rect 1630 -3575 1750 -3570
rect 1630 -3720 1750 -3710
rect 1630 -3755 1710 -3720
rect 1745 -3755 1750 -3720
rect 1630 -3760 1750 -3755
rect 1630 -3905 1750 -3895
rect 1630 -3940 1710 -3905
rect 1745 -3940 1750 -3905
rect 1630 -3945 1750 -3940
rect 1630 -4090 1750 -4080
rect 1630 -4125 1710 -4090
rect 1745 -4125 1750 -4090
rect 1630 -4130 1750 -4125
rect 1630 -4275 1750 -4265
rect 1630 -4310 1710 -4275
rect 1745 -4310 1750 -4275
rect 1630 -4315 1750 -4310
<< end >>
